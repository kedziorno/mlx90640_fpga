----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:12:21 02/09/2023 
-- Design Name: 
-- Module Name:    mem_unsigned1024 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
----library UNISIM;
----use UNISIM.VComponents.all;

entity mem_unsigned1024 is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_value : in std_logic_vector (9 downto 0); -- input hex from 0 to 1024
o_value : out std_logic_vector (31 downto 0) -- output signed 0 to 1024 in SP float
);
end mem_unsigned1024;

architecture Behavioral of mem_unsigned1024 is

COMPONENT mem_ramb16_s36_x2
generic (
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0a : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0b : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0c : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0d : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0e : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0f : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
);
PORT(
DO : OUT  std_logic_vector(31 downto 0);
DOP : OUT  std_logic_vector(3 downto 0);
ADDR : IN  std_logic_vector(9 downto 0);
CLK : IN  std_logic;
DI : IN  std_logic_vector(31 downto 0);
DIP : IN  std_logic_vector(3 downto 0);
EN : IN  std_logic;
SSR : IN  std_logic;
WE : IN  std_logic
);
END COMPONENT mem_ramb16_s36_x2;

begin

inst_unsigned1024 : mem_ramb16_s36_x2 
GENERIC MAP (
INIT_00 => X"40e0000040c0000040a000004080000040400000400000003f80000000000000",       
INIT_01 => X"4170000041600000415000004140000041300000412000004110000041000000",
INIT_02 => X"41b8000041b0000041a8000041a0000041980000419000004188000041800000",
INIT_03 => X"41f8000041f0000041e8000041e0000041d8000041d0000041c8000041c00000",
INIT_04 => X"421c0000421800004214000042100000420c0000420800004204000042000000",
INIT_05 => X"423c0000423800004234000042300000422c0000422800004224000042200000",
INIT_06 => X"425c0000425800004254000042500000424c0000424800004244000042400000",
INIT_07 => X"427c0000427800004274000042700000426c0000426800004264000042600000",
INIT_08 => X"428e0000428c0000428a00004288000042860000428400004282000042800000",
INIT_09 => X"429e0000429c0000429a00004298000042960000429400004292000042900000",
INIT_0a => X"42ae000042ac000042aa000042a8000042a6000042a4000042a2000042a00000",
INIT_0b => X"42be000042bc000042ba000042b8000042b6000042b4000042b2000042b00000",
INIT_0c => X"42ce000042cc000042ca000042c8000042c6000042c4000042c2000042c00000",
INIT_0d => X"42de000042dc000042da000042d8000042d6000042d4000042d2000042d00000",
INIT_0e => X"42ee000042ec000042ea000042e8000042e6000042e4000042e2000042e00000",
INIT_0f => X"42fe000042fc000042fa000042f8000042f6000042f4000042f2000042f00000",
INIT_10 => X"4307000043060000430500004304000043030000430200004301000043000000",
INIT_11 => X"430f0000430e0000430d0000430c0000430b0000430a00004309000043080000",
INIT_12 => X"4317000043160000431500004314000043130000431200004311000043100000",
INIT_13 => X"431f0000431e0000431d0000431c0000431b0000431a00004319000043180000",
INIT_14 => X"4327000043260000432500004324000043230000432200004321000043200000",
INIT_15 => X"432f0000432e0000432d0000432c0000432b0000432a00004329000043280000",
INIT_16 => X"4337000043360000433500004334000043330000433200004331000043300000",
INIT_17 => X"433f0000433e0000433d0000433c0000433b0000433a00004339000043380000",
INIT_18 => X"4347000043460000434500004344000043430000434200004341000043400000",
INIT_19 => X"434f0000434e0000434d0000434c0000434b0000434a00004349000043480000",
INIT_1a => X"4357000043560000435500004354000043530000435200004351000043500000",
INIT_1b => X"435f0000435e0000435d0000435c0000435b0000435a00004359000043580000",
INIT_1c => X"4367000043660000436500004364000043630000436200004361000043600000",
INIT_1d => X"436f0000436e0000436d0000436c0000436b0000436a00004369000043680000",
INIT_1e => X"4377000043760000437500004374000043730000437200004371000043700000",
INIT_1f => X"437f0000437e0000437d0000437c0000437b0000437a00004379000043780000",
INIT_20 => X"4383800043830000438280004382000043818000438100004380800043800000",
INIT_21 => X"4387800043870000438680004386000043858000438500004384800043840000",
INIT_22 => X"438b8000438b0000438a8000438a000043898000438900004388800043880000",
INIT_23 => X"438f8000438f0000438e8000438e0000438d8000438d0000438c8000438c0000",
INIT_24 => X"4393800043930000439280004392000043918000439100004390800043900000",
INIT_25 => X"4397800043970000439680004396000043958000439500004394800043940000",
INIT_26 => X"439b8000439b0000439a8000439a000043998000439900004398800043980000",
INIT_27 => X"439f8000439f0000439e8000439e0000439d8000439d0000439c8000439c0000",
INIT_28 => X"43a3800043a3000043a2800043a2000043a1800043a1000043a0800043a00000",
INIT_29 => X"43a7800043a7000043a6800043a6000043a5800043a5000043a4800043a40000",
INIT_2a => X"43ab800043ab000043aa800043aa000043a9800043a9000043a8800043a80000",
INIT_2b => X"43af800043af000043ae800043ae000043ad800043ad000043ac800043ac0000",
INIT_2c => X"43b3800043b3000043b2800043b2000043b1800043b1000043b0800043b00000",
INIT_2d => X"43b7800043b7000043b6800043b6000043b5800043b5000043b4800043b40000",
INIT_2e => X"43bb800043bb000043ba800043ba000043b9800043b9000043b8800043b80000",
INIT_2f => X"43bf800043bf000043be800043be000043bd800043bd000043bc800043bc0000",
INIT_30 => X"43c3800043c3000043c2800043c2000043c1800043c1000043c0800043c00000",
INIT_31 => X"43c7800043c7000043c6800043c6000043c5800043c5000043c4800043c40000",
INIT_32 => X"43cb800043cb000043ca800043ca000043c9800043c9000043c8800043c80000",
INIT_33 => X"43cf800043cf000043ce800043ce000043cd800043cd000043cc800043cc0000",
INIT_34 => X"43d3800043d3000043d2800043d2000043d1800043d1000043d0800043d00000",
INIT_35 => X"43d7800043d7000043d6800043d6000043d5800043d5000043d4800043d40000",
INIT_36 => X"43db800043db000043da800043da000043d9800043d9000043d8800043d80000",
INIT_37 => X"43df800043df000043de800043de000043dd800043dd000043dc800043dc0000",
INIT_38 => X"43e3800043e3000043e2800043e2000043e1800043e1000043e0800043e00000",
INIT_39 => X"43e7800043e7000043e6800043e6000043e5800043e5000043e4800043e40000",
INIT_3a => X"43eb800043eb000043ea800043ea000043e9800043e9000043e8800043e80000",
INIT_3b => X"43ef800043ef000043ee800043ee000043ed800043ed000043ec800043ec0000",
INIT_3c => X"43f3800043f3000043f2800043f2000043f1800043f1000043f0800043f00000",
INIT_3d => X"43f7800043f7000043f6800043f6000043f5800043f5000043f4800043f40000",
INIT_3e => X"43fb800043fb000043fa800043fa000043f9800043f9000043f8800043f80000",
INIT_3f => X"43ff800043ff000043fe800043fe000043fd800043fd000043fc800043fc0000",
INIT_40 => X"4401c0004401800044014000440100004400c000440080004400400044000000",
INIT_41 => X"4403c0004403800044034000440300004402c000440280004402400044020000",
INIT_42 => X"4405c0004405800044054000440500004404c000440480004404400044040000",
INIT_43 => X"4407c0004407800044074000440700004406c000440680004406400044060000",
INIT_44 => X"4409c0004409800044094000440900004408c000440880004408400044080000",
INIT_45 => X"440bc000440b8000440b4000440b0000440ac000440a8000440a4000440a0000",
INIT_46 => X"440dc000440d8000440d4000440d0000440cc000440c8000440c4000440c0000",
INIT_47 => X"440fc000440f8000440f4000440f0000440ec000440e8000440e4000440e0000",
INIT_48 => X"4411c0004411800044114000441100004410c000441080004410400044100000",
INIT_49 => X"4413c0004413800044134000441300004412c000441280004412400044120000",
INIT_4a => X"4415c0004415800044154000441500004414c000441480004414400044140000",
INIT_4b => X"4417c0004417800044174000441700004416c000441680004416400044160000",
INIT_4c => X"4419c0004419800044194000441900004418c000441880004418400044180000",
INIT_4d => X"441bc000441b8000441b4000441b0000441ac000441a8000441a4000441a0000",
INIT_4e => X"441dc000441d8000441d4000441d0000441cc000441c8000441c4000441c0000",
INIT_4f => X"441fc000441f8000441f4000441f0000441ec000441e8000441e4000441e0000",
INIT_50 => X"4421c0004421800044214000442100004420c000442080004420400044200000",
INIT_51 => X"4423c0004423800044234000442300004422c000442280004422400044220000",
INIT_52 => X"4425c0004425800044254000442500004424c000442480004424400044240000",
INIT_53 => X"4427c0004427800044274000442700004426c000442680004426400044260000",
INIT_54 => X"4429c0004429800044294000442900004428c000442880004428400044280000",
INIT_55 => X"442bc000442b8000442b4000442b0000442ac000442a8000442a4000442a0000",
INIT_56 => X"442dc000442d8000442d4000442d0000442cc000442c8000442c4000442c0000",
INIT_57 => X"442fc000442f8000442f4000442f0000442ec000442e8000442e4000442e0000",
INIT_58 => X"4431c0004431800044314000443100004430c000443080004430400044300000",
INIT_59 => X"4433c0004433800044334000443300004432c000443280004432400044320000",
INIT_5a => X"4435c0004435800044354000443500004434c000443480004434400044340000",
INIT_5b => X"4437c0004437800044374000443700004436c000443680004436400044360000",
INIT_5c => X"4439c0004439800044394000443900004438c000443880004438400044380000",
INIT_5d => X"443bc000443b8000443b4000443b0000443ac000443a8000443a4000443a0000",
INIT_5e => X"443dc000443d8000443d4000443d0000443cc000443c8000443c4000443c0000",
INIT_5f => X"443fc000443f8000443f4000443f0000443ec000443e8000443e4000443e0000",
INIT_60 => X"4441c0004441800044414000444100004440c000444080004440400044400000",
INIT_61 => X"4443c0004443800044434000444300004442c000444280004442400044420000",
INIT_62 => X"4445c0004445800044454000444500004444c000444480004444400044440000",
INIT_63 => X"4447c0004447800044474000444700004446c000444680004446400044460000",
INIT_64 => X"4449c0004449800044494000444900004448c000444880004448400044480000",
INIT_65 => X"444bc000444b8000444b4000444b0000444ac000444a8000444a4000444a0000",
INIT_66 => X"444dc000444d8000444d4000444d0000444cc000444c8000444c4000444c0000",
INIT_67 => X"444fc000444f8000444f4000444f0000444ec000444e8000444e4000444e0000",
INIT_68 => X"4451c0004451800044514000445100004450c000445080004450400044500000",
INIT_69 => X"4453c0004453800044534000445300004452c000445280004452400044520000",
INIT_6a => X"4455c0004455800044554000445500004454c000445480004454400044540000",
INIT_6b => X"4457c0004457800044574000445700004456c000445680004456400044560000",
INIT_6c => X"4459c0004459800044594000445900004458c000445880004458400044580000",
INIT_6d => X"445bc000445b8000445b4000445b0000445ac000445a8000445a4000445a0000",
INIT_6e => X"445dc000445d8000445d4000445d0000445cc000445c8000445c4000445c0000",
INIT_6f => X"445fc000445f8000445f4000445f0000445ec000445e8000445e4000445e0000",
INIT_70 => X"4461c0004461800044614000446100004460c000446080004460400044600000",
INIT_71 => X"4463c0004463800044634000446300004462c000446280004462400044620000",
INIT_72 => X"4465c0004465800044654000446500004464c000446480004464400044640000",
INIT_73 => X"4467c0004467800044674000446700004466c000446680004466400044660000",
INIT_74 => X"4469c0004469800044694000446900004468c000446880004468400044680000",
INIT_75 => X"446bc000446b8000446b4000446b0000446ac000446a8000446a4000446a0000",
INIT_76 => X"446dc000446d8000446d4000446d0000446cc000446c8000446c4000446c0000",
INIT_77 => X"446fc000446f8000446f4000446f0000446ec000446e8000446e4000446e0000",
INIT_78 => X"4471c0004471800044714000447100004470c000447080004470400044700000",
INIT_79 => X"4473c0004473800044734000447300004472c000447280004472400044720000",
INIT_7a => X"4475c0004475800044754000447500004474c000447480004474400044740000",
INIT_7b => X"4477c0004477800044774000447700004476c000447680004476400044760000",
INIT_7c => X"4479c0004479800044794000447900004478c000447880004478400044780000",
INIT_7d => X"447bc000447b8000447b4000447b0000447ac000447a8000447a4000447a0000",
INIT_7e => X"447dc000447d8000447d4000447d0000447cc000447c8000447c4000447c0000",
INIT_7f => X"447fc000447f8000447f4000447f0000447ec000447e8000447e4000447e0000"
)
PORT MAP (
DO => o_value,
DOP => open,
ADDR => i_value,
CLK => i_clock,
DI => (others => '0'),
DIP => (others => '0'),
EN => '1',
SSR => i_reset,
WE => '0'
);

end Behavioral;

