----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:44:29 02/05/2023 
-- Design Name: 
-- Module Name:    mem_signedFF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mem_signedFF is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_value : in std_logic_vector (7 downto 0); -- input hex from 0 to 255
o_value : out std_logic_vector (31 downto 0) -- output signed -128 to 127 in SP float
);
end mem_signedFF;

architecture Behavioral of mem_signedFF is

begin

inst_mem_signedFF : RAMB16_S36
generic map (
INIT => X"0", -- Value of output RAM registers at startup
SRVAL => X"0", -- Output value upon SSR assertion
WRITE_MODE => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
-- The following INIT_xx declarations specify the intial contents of the RAM
-- Address 0 to 4095
INIT_00 => X"40e0000040c0000040a000004080000040400000400000003f80000000000000",
INIT_01 => X"4170000041600000415000004140000041300000412000004110000041000000",
INIT_02 => X"41b8000041b0000041a8000041a0000041980000419000004188000041800000",
INIT_03 => X"41f8000041f0000041e8000041e0000041d8000041d0000041c8000041c00000",
INIT_04 => X"421c0000421800004214000042100000420c0000420800004204000042000000",
INIT_05 => X"423c0000423800004234000042300000422c0000422800004224000042200000",
INIT_06 => X"425c0000425800004254000042500000424c0000424800004244000042400000",
INIT_07 => X"427c0000427800004274000042700000426c0000426800004264000042600000",
INIT_08 => X"428e0000428c0000428a00004288000042860000428400004282000042800000",
INIT_09 => X"429e0000429c0000429a00004298000042960000429400004292000042900000",
INIT_0a => X"42ae000042ac000042aa000042a8000042a6000042a4000042a2000042a00000",
INIT_0b => X"42be000042bc000042ba000042b8000042b6000042b4000042b2000042b00000",
INIT_0c => X"42ce000042cc000042ca000042c8000042c6000042c4000042c2000042c00000",
INIT_0d => X"42de000042dc000042da000042d8000042d6000042d4000042d2000042d00000",
INIT_0e => X"42ee000042ec000042ea000042e8000042e6000042e4000042e2000042e00000",
INIT_0f => X"42fe000042fc000042fa000042f8000042f6000042f4000042f2000042f00000",
INIT_10 => X"c2f20000c2f40000c2f60000c2f80000c2fa0000c2fc0000c2fe0000c3000000",
INIT_11 => X"c2e20000c2e40000c2e60000c2e80000c2ea0000c2ec0000c2ee0000c2f00000",
INIT_12 => X"c2d20000c2d40000c2d60000c2d80000c2da0000c2dc0000c2de0000c2e00000",
INIT_13 => X"c2c20000c2c40000c2c60000c2c80000c2ca0000c2cc0000c2ce0000c2d00000",
INIT_14 => X"c2b20000c2b40000c2b60000c2b80000c2ba0000c2bc0000c2be0000c2c00000",
INIT_15 => X"c2a20000c2a40000c2a60000c2a80000c2aa0000c2ac0000c2ae0000c2b00000",
INIT_16 => X"c2920000c2940000c2960000c2980000c29a0000c29c0000c29e0000c2a00000",
INIT_17 => X"c2820000c2840000c2860000c2880000c28a0000c28c0000c28e0000c2900000",
INIT_18 => X"c2640000c2680000c26c0000c2700000c2740000c2780000c27c0000c2800000",
INIT_19 => X"c2440000c2480000c24c0000c2500000c2540000c2580000c25c0000c2600000",
INIT_1a => X"c2240000c2280000c22c0000c2300000c2340000c2380000c23c0000c2400000",
INIT_1b => X"c2040000c2080000c20c0000c2100000c2140000c2180000c21c0000c2200000",
INIT_1c => X"c1c80000c1d00000c1d80000c1e00000c1e80000c1f00000c1f80000c2000000",
INIT_1d => X"c1880000c1900000c1980000c1a00000c1a80000c1b00000c1b80000c1c00000",
INIT_1e => X"c1100000c1200000c1300000c1400000c1500000c1600000c1700000c1800000",
INIT_1f => X"bf800000c0000000c0400000c0800000c0a00000c0c00000c0e00000c1000000",
-- Address 8192 to 12287
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 12288 to 16383
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
DO => o_value, -- 1-bit Data Output
DOP => open, -- 1-bit Data Output
ADDR => "0"&i_value, -- 14-bit Address Input
CLK => i_clock, -- Clock
DI => (others => '0'), -- 1-bit Data Input
DIP => (others => '0'), -- 1-bit Data Input
EN => '1', -- RAM Enable Input
SSR => i_reset, -- Synchronous Set/Reset Input
WE => '0' -- Write Enable Input
);
-- End of RAMB16_S1_inst instantiation

end Behavioral;

