idle,5

address,33,1
data,ff,0
data,ff,0
data,ff,0
data,ff,0

idle,1

address,33,0
data,ff,0
data,ff,0

idle,3

address,33,0
data,ff,0
data,ff,1

idle,17

idle,15

address,33,0
data,ff,0
data,54,1
data,ab,0
data,2a,1
data,d5,0
data,00,1
data,ff,0

idle,11

address,33,1
data,ff,1
data,32,1
data,cd,1
data,54,1
data,ab,1
data,2a,1

idle,13

address,33,1
data,ff,0
data,00,0
data,d5,0
data,2a,1
data,ab,0
data,54,0
data,00,0
data,ff,1

idle,13

