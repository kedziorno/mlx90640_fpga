
package p_fphdl_package3 is


end p_fphdl_package3;

package body p_fphdl_package3 is


end p_fphdl_package3;
