----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:20:04 12/23/2022 
-- Design Name: 
-- Module Name:    mem_kvptat_ktptat - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mem_kvptat_ktptat is
port (
	i_clock : in std_logic;
	i_reset : in std_logic;
	i_address : in std_logic_vector(14 downto 0);
	o_data_kvptat : out std_logic_vector(31 downto 0);
	o_data_ktptat : out std_logic_vector(31 downto 0)
);
end mem_kvptat_ktptat;

architecture Behavioral of mem_kvptat_ktptat is

component RAMB16 is
generic (
DOA_REG : integer := 0 ;
DOB_REG : integer := 0 ;
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_A : bit_vector := X"000000000";
INIT_B : bit_vector := X"000000000";
INIT_FILE : string := "NONE";
INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INVERT_CLK_DOA_REG : boolean := false;
INVERT_CLK_DOB_REG : boolean := false;
RAM_EXTENSION_A : string := "NONE";
RAM_EXTENSION_B : string := "NONE";
READ_WIDTH_A : integer := 0;
READ_WIDTH_B : integer := 0;
SIM_COLLISION_CHECK : string := "ALL";
SRVAL_A  : bit_vector := X"000000000";
SRVAL_B  : bit_vector := X"000000000";
WRITE_MODE_A : string := "WRITE_FIRST";
WRITE_MODE_B : string := "WRITE_FIRST";
WRITE_WIDTH_A : integer := 0;
WRITE_WIDTH_B : integer := 0
);
port(
CASCADEOUTA  : out  std_ulogic;
CASCADEOUTB  : out  std_ulogic;
DOA          : out std_logic_vector (31 downto 0);
DOB          : out std_logic_vector (31 downto 0);
DOPA         : out std_logic_vector (3 downto 0);
DOPB         : out std_logic_vector (3 downto 0);
ADDRA        : in  std_logic_vector (14 downto 0);
ADDRB        : in  std_logic_vector (14 downto 0);
CASCADEINA   : in  std_ulogic;
CASCADEINB   : in  std_ulogic;
CLKA         : in  std_ulogic;
CLKB         : in  std_ulogic;
DIA          : in  std_logic_vector (31 downto 0);
DIB          : in  std_logic_vector (31 downto 0);
DIPA         : in  std_logic_vector (3 downto 0);
DIPB         : in  std_logic_vector (3 downto 0);
ENA          : in  std_ulogic;
ENB          : in  std_ulogic;
REGCEA       : in  std_ulogic;
REGCEB       : in  std_ulogic;
SSRA         : in  std_ulogic;
SSRB         : in  std_ulogic;
WEA          : in  std_logic_vector (3 downto 0);
WEB          : in  std_logic_vector (3 downto 0)
);
end component RAMB16;

signal odata_kvptat : std_logic_vector(31 downto 0);
signal odata_ktptat : std_logic_vector(31 downto 0);
signal address_kvptat : std_logic_vector(14 downto 0);
signal address_ktptat : std_logic_vector(14 downto 0);

begin

--p0 : process (i_address) is
--begin
--	address_kvptat <= std_logic_vector(to_unsigned(to_integer(unsigned(i_address)) * 32,15));
--end process p0;

p1 : process (i_address) is
begin
	address_ktptat <= std_logic_vector(to_unsigned(((to_integer(unsigned(i_address))) * 16),15));
end process p1;

o_data_kvptat <= odata_kvptat;
o_data_ktptat <= odata_ktptat(15 downto 0) & x"0000";

inst_mem_kvdd : RAMB16
generic map (
DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
INIT_A => X"000000000", -- Initial values on A output port
INIT_B => X"000000000", -- Initial values on B output port
INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
READ_WIDTH_A => 36, -- Valid values are 1,2,4,9,18 or 36
READ_WIDTH_B => 36, -- Valid values are 1,2,4,9,18 or 36
SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
WRITE_MODE_A => "NO_CHANGE", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_MODE_B => "NO_CHANGE", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_WIDTH_A => 36, -- Valid values are 1,2,4,9,18 or 36
WRITE_WIDTH_B => 36, -- Valid values are 1,2,4,9,18 or 36

-- page36 11.2.2.3
-- ktptat 0x0-0x3FF
INIT_00 => X"3f803f003e803e003d803d003c803c003b003a00390038003600340030000000",   
INIT_01 => X"43c043804340430042c042804240420041c041804140410040c0408040404000",
INIT_02 => X"45e045c045a04580456045404520450044e044c044a044804460444044204400",
INIT_03 => X"47e047c047a04780476047404720470046e046c046a046804660464046204600",
INIT_04 => X"48f048e048d048c048b048a04890488048704860485048404830482048104800",
INIT_05 => X"49f049e049d049c049b049a04990498049704960495049404930492049104900",
INIT_06 => X"4af04ae04ad04ac04ab04aa04a904a804a704a604a504a404a304a204a104a00",
INIT_07 => X"4bf04be04bd04bc04bb04ba04b904b804b704b604b504b404b304b204b104b00",
INIT_08 => X"4c784c704c684c604c584c504c484c404c384c304c284c204c184c104c084c00",
INIT_09 => X"4cf84cf04ce84ce04cd84cd04cc84cc04cb84cb04ca84ca04c984c904c884c80",
INIT_0a => X"4d784d704d684d604d584d504d484d404d384d304d284d204d184d104d084d00",
INIT_0b => X"4df84df04de84de04dd84dd04dc84dc04db84db04da84da04d984d904d884d80",
INIT_0c => X"4e784e704e684e604e584e504e484e404e384e304e284e204e184e104e084e00",
INIT_0d => X"4ef84ef04ee84ee04ed84ed04ec84ec04eb84eb04ea84ea04e984e904e884e80",
INIT_0e => X"4f784f704f684f604f584f504f484f404f384f304f284f204f184f104f084f00",
INIT_0f => X"4ff84ff04fe84fe04fd84fd04fc84fc04fb84fb04fa84fa04f984f904f884f80",
INIT_10 => X"503c503850345030502c502850245020501c501850145010500c500850045000",
INIT_11 => X"507c507850745070506c506850645060505c505850545050504c504850445040",
INIT_12 => X"50bc50b850b450b050ac50a850a450a0509c509850945090508c508850845080",
INIT_13 => X"50fc50f850f450f050ec50e850e450e050dc50d850d450d050cc50c850c450c0",
INIT_14 => X"513c513851345130512c512851245120511c511851145110510c510851045100",
INIT_15 => X"517c517851745170516c516851645160515c515851545150514c514851445140",
INIT_16 => X"51bc51b851b451b051ac51a851a451a0519c519851945190518c518851845180",
INIT_17 => X"51fc51f851f451f051ec51e851e451e051dc51d851d451d051cc51c851c451c0",
INIT_18 => X"523c523852345230522c522852245220521c521852145210520c520852045200",
INIT_19 => X"527c527852745270526c526852645260525c525852545250524c524852445240",
INIT_1a => X"52bc52b852b452b052ac52a852a452a0529c529852945290528c528852845280",
INIT_1b => X"52fc52f852f452f052ec52e852e452e052dc52d852d452d052cc52c852c452c0",
INIT_1c => X"533c533853345330532c532853245320531c531853145310530c530853045300",
INIT_1d => X"537c537853745370536c536853645360535c535853545350534c534853445340",
INIT_1e => X"53bc53b853b453b053ac53a853a453a0539c539853945390538c538853845380",
INIT_1f => X"53fc53f853f453f053ec53e853e453e053dc53d853d453d053cc53c853c453c0",
INIT_20 => X"d3c4d3c8d3ccd3d0d3d4d3d8d3dcd3e0d3e4d3e8d3ecd3f0d3f4d3f8d3fcd400",
INIT_21 => X"d384d388d38cd390d394d398d39cd3a0d3a4d3a8d3acd3b0d3b4d3b8d3bcd3c0",
INIT_22 => X"d344d348d34cd350d354d358d35cd360d364d368d36cd370d374d378d37cd380",
INIT_23 => X"d304d308d30cd310d314d318d31cd320d324d328d32cd330d334d338d33cd340",
INIT_24 => X"d2c4d2c8d2ccd2d0d2d4d2d8d2dcd2e0d2e4d2e8d2ecd2f0d2f4d2f8d2fcd300",
INIT_25 => X"d284d288d28cd290d294d298d29cd2a0d2a4d2a8d2acd2b0d2b4d2b8d2bcd2c0",
INIT_26 => X"d244d248d24cd250d254d258d25cd260d264d268d26cd270d274d278d27cd280",
INIT_27 => X"d204d208d20cd210d214d218d21cd220d224d228d22cd230d234d238d23cd240",
INIT_28 => X"d1c4d1c8d1ccd1d0d1d4d1d8d1dcd1e0d1e4d1e8d1ecd1f0d1f4d1f8d1fcd200",
INIT_29 => X"d184d188d18cd190d194d198d19cd1a0d1a4d1a8d1acd1b0d1b4d1b8d1bcd1c0",
INIT_2a => X"d144d148d14cd150d154d158d15cd160d164d168d16cd170d174d178d17cd180",
INIT_2b => X"d104d108d10cd110d114d118d11cd120d124d128d12cd130d134d138d13cd140",
INIT_2c => X"d0c4d0c8d0ccd0d0d0d4d0d8d0dcd0e0d0e4d0e8d0ecd0f0d0f4d0f8d0fcd100",
INIT_2d => X"d084d088d08cd090d094d098d09cd0a0d0a4d0a8d0acd0b0d0b4d0b8d0bcd0c0",
INIT_2e => X"d044d048d04cd050d054d058d05cd060d064d068d06cd070d074d078d07cd080",
INIT_2f => X"d004d008d00cd010d014d018d01cd020d024d028d02cd030d034d038d03cd040",
INIT_30 => X"cf88cf90cf98cfa0cfa8cfb0cfb8cfc0cfc8cfd0cfd8cfe0cfe8cff0cff8d000",
INIT_31 => X"cf08cf10cf18cf20cf28cf30cf38cf40cf48cf50cf58cf60cf68cf70cf78cf80",
INIT_32 => X"ce88ce90ce98cea0cea8ceb0ceb8cec0cec8ced0ced8cee0cee8cef0cef8cf00",
INIT_33 => X"ce08ce10ce18ce20ce28ce30ce38ce40ce48ce50ce58ce60ce68ce70ce78ce80",
INIT_34 => X"cd88cd90cd98cda0cda8cdb0cdb8cdc0cdc8cdd0cdd8cde0cde8cdf0cdf8ce00",
INIT_35 => X"cd08cd10cd18cd20cd28cd30cd38cd40cd48cd50cd58cd60cd68cd70cd78cd80",
INIT_36 => X"cc88cc90cc98cca0cca8ccb0ccb8ccc0ccc8ccd0ccd8cce0cce8ccf0ccf8cd00",
INIT_37 => X"cc08cc10cc18cc20cc28cc30cc38cc40cc48cc50cc58cc60cc68cc70cc78cc80",
INIT_38 => X"cb10cb20cb30cb40cb50cb60cb70cb80cb90cba0cbb0cbc0cbd0cbe0cbf0cc00",
INIT_39 => X"ca10ca20ca30ca40ca50ca60ca70ca80ca90caa0cab0cac0cad0cae0caf0cb00",
INIT_3a => X"c910c920c930c940c950c960c970c980c990c9a0c9b0c9c0c9d0c9e0c9f0ca00",
INIT_3b => X"c810c820c830c840c850c860c870c880c890c8a0c8b0c8c0c8d0c8e0c8f0c900",
INIT_3c => X"c620c640c660c680c6a0c6c0c6e0c700c720c740c760c780c7a0c7c0c7e0c800",
INIT_3d => X"c420c440c460c480c4a0c4c0c4e0c500c520c540c560c580c5a0c5c0c5e0c600",
INIT_3e => X"c040c080c0c0c100c140c180c1c0c200c240c280c2c0c300c340c380c3c0c400",
INIT_3f => X"b000b400b600b800b900ba00bb00bc00bc80bd00bd80be00be80bf00bf80c000",
INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
)
port map (
CASCADEOUTA => open, -- 1-bit cascade output
CASCADEOUTB => open, -- 1-bit cascade output
DOA => odata_kvptat, -- 32-bit A port Data Output
DOB => odata_ktptat, -- 32-bit B port Data Output
DOPA => open, -- 4-bit A port Parity Output
DOPB => open, -- 4-bit B port Parity Output
ADDRA => address_kvptat, -- 15-bit A port Address Input
ADDRB => address_ktptat, -- 15-bit B port Address Input
CASCADEINA => '0', -- 1-bit cascade A input
CASCADEINB => '0', -- 1-bit cascade B input
CLKA => i_clock, -- Port A Clock
CLKB => i_clock, -- Port B Clock
DIA => (others => '0'), -- 32-bit A port Data Input
DIB => (others => '0'), -- 32-bit B port Data Input
DIPA => (others => '0'), -- 4-bit A port parity Input
DIPB => (others => '0'), -- 4-bit B port parity Input
ENA => '1', -- 1-bit A port Enable Input
ENB => '1', -- 1-bit B port Enable Input
REGCEA => '1', -- 1-bit A port register enable input
REGCEB => '1', -- 1-bit B port register enable input
SSRA => i_reset, -- 1-bit A port Synchronous Set/Reset Input
SSRB => i_reset, -- 1-bit B port Synchronous Set/Reset Input
WEA => (others => '0'), -- 4-bit A port Write Enable Input
WEB => (others => '0') -- 4-bit B port Write Enable Input
);

--RAMB16
--generic map (
--DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
--DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
--INIT_A => X"000000000", -- Initial values on A output port
--INIT_B => X"000000000", -- Initial values on B output port
--INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
--INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
--RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--READ_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36
--READ_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
--SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
--SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
--WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
--WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
--WRITE_WIDTH_A => 2, -- Valid values are 1,2,4,9,18 or 36
--WRITE_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
--INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
--)
--port map (
--CASCADEOUTA => CASCADEOUTA, -- 1-bit cascade output
--CASCADEOUTB => CASCADEOUTB, -- 1-bit cascade output
--DOA => DOA, -- 32-bit A port Data Output
--DOB => DOB, -- 32-bit B port Data Output
--DOPA => DOPA, -- 4-bit A port Parity Output
--DOPB => DOPB, -- 4-bit B port Parity Output
--ADDRA => ADDRA, -- 15-bit A port Address Input
--ADDRB => ADDRB, -- 15-bit B port Address Input
--CASCADEINA => CASCADEINA, -- 1-bit cascade A input
--CASCADEINB => CASCADEINB, -- 1-bit cascade B input
--CLKA => CLKA, -- Port A Clock
--CLKB => CLKB, -- Port B Clock
--DIA => DIA, -- 32-bit A port Data Input
--DIB => DIB, -- 32-bit B port Data Input
--DIPA => DIPA, -- 4-bit A port parity Input
--DIPB => DIPB, -- 4-bit B port parity Input
--ENA => ENA, -- 1-bit A port Enable Input
--ENB => ENB, -- 1-bit B port Enable Input
--REGCEA => REGCEA, -- 1-bit A port register enable input
--REGCEB => REGCEB, -- 1-bit B port register enable input
--SSRA => SSRA, -- 1-bit A port Synchronous Set/Reset Input
--SSRB => SSRB, -- 1-bit B port Synchronous Set/Reset Input
--WEA => WEA, -- 4-bit A port Write Enable Input
--WEB => WEB -- 4-bit B port Write Enable Input
--);

end Behavioral;
