library IEEE;
use IEEE.STD_LOGIC_1164.all;

package colormap_pkg is

type rom_type is array (-128 to 127) of std_logic_vector (23 downto 0);
constant colormap_rom : rom_type := (
x"04001f",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"04001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"05001e",
x"06001e",
x"06001e",
x"06001e",
x"06001e",
x"06001e",
x"06001e",
x"06001e",
x"06001e",
x"06001d",
x"06001d",
x"06001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"07001d",
x"08001d",
x"08001c",
x"08001c",
x"08001c",
x"08001c",
x"08001c",
x"08001c",
x"08001c",
x"08001c",
x"09001c",
x"09001c",
x"09001c",
x"09001b",
x"09001b",
x"09001b",
x"09001b",
x"09001b",
x"09001b",
x"0a001b",
x"0a001b",
x"0a001b",
x"0a001b",
x"0a001a",
x"0a001a",
x"0a001a",
x"0a001a",
x"0b001a",
x"0b001a",
x"0b001a",
x"0b001a",
x"0b0019",
x"0b0019",
x"0b0019",
x"0b0019",
x"0c0019",
x"0c0019",
x"0c0019",
x"0c0019",
x"0c0018",
x"0c0018",
x"0c0018",
x"0c0018",
x"0d0018",
x"0d0018",
x"0d0018",
x"0d0018",
x"0d0017",
x"0d0017",
x"0d0017",
x"0e0017",
x"0e0017",
x"0e0017",
x"0e0017",
x"0e0016",
x"0e0016",
x"0e0016",
x"0f0016",
x"0f0016",
x"0f0016",
x"0f0016",
x"0f0016",
x"0f0015",
x"0f0015",
x"100015",
x"100015",
x"100015",
x"100015",
x"100014",
x"100014",
x"100014",
x"110014",
x"110014",
x"110014",
x"110014",
x"110013",
x"110013",
x"110013",
x"120013",
x"120013",
x"120013",
x"120013",
x"120012",
x"120012",
x"120012",
x"130012",
x"130012",
x"130012",
x"130012",
x"130011",
x"130011",
x"130011",
x"140011",
x"140011",
x"140011",
x"140011",
x"140010",
x"140010",
x"140010",
x"150010",
x"150010",
x"150010",
x"150010",
x"15000f",
x"15000f",
x"16000f",
x"16000f",
x"16000f",
x"16000f",
x"16000f",
x"16000e",
x"16000e",
x"16000e",
x"17000e",
x"17000e",
x"17000e",
x"17000e",
x"17000d",
x"17000d",
x"17000d",
x"18000d",
x"18000d",
x"18000d",
x"18000d",
x"18000c",
x"18000c",
x"18000c",
x"18000c",
x"19000c",
x"19000c",
x"19000c",
x"19000c",
x"19000b",
x"19000b",
x"19000b",
x"19000b",
x"1a000b",
x"1a000b",
x"1a000b",
x"1a000b",
x"1a000a",
x"1a000a",
x"1a000a",
x"1a000a",
x"1b000a",
x"1b000a",
x"1b000a",
x"1b000a",
x"1b0009",
x"1b0009",
x"1b0009",
x"1b0009",
x"1b0009",
x"1b0009",
x"1c0009",
x"1c0009",
x"1c0009",
x"1c0008",
x"1c0008",
x"1c0008",
x"1c0008",
x"1c0008",
x"1c0008",
x"1c0008",
x"1c0008",
x"1d0008",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0007",
x"1d0006",
x"1d0006",
x"1d0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0006",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0005",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004",
x"1e0004"
);

end colormap_pkg;

package body colormap_pkg is
 
end colormap_pkg;
