----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:03:24 12/13/2022 
-- Design Name: 
-- Module Name:    mem_kvdd_vdd25 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mem_kvdd_vdd25 is
port (
	i_clock : in std_logic;
	i_reset : in std_logic;
	i_address : in std_logic_vector(7 downto 0);
	o_data_kvdd : out std_logic_vector(15 downto 0);
	o_data_vdd25 : out std_logic_vector(15 downto 0)
);
end entity mem_kvdd_vdd25;

architecture Behavioral of mem_kvdd_vdd25 is

component RAMB16 is
generic (
DOA_REG : integer := 0 ;
DOB_REG : integer := 0 ;
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_A : bit_vector := X"000000000";
INIT_B : bit_vector := X"000000000";
INIT_FILE : string := "NONE";
INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INVERT_CLK_DOA_REG : boolean := false;
INVERT_CLK_DOB_REG : boolean := false;
RAM_EXTENSION_A : string := "NONE";
RAM_EXTENSION_B : string := "NONE";
READ_WIDTH_A : integer := 0;
READ_WIDTH_B : integer := 0;
SIM_COLLISION_CHECK : string := "ALL";
SRVAL_A  : bit_vector := X"000000000";
SRVAL_B  : bit_vector := X"000000000";
WRITE_MODE_A : string := "WRITE_FIRST";
WRITE_MODE_B : string := "WRITE_FIRST";
WRITE_WIDTH_A : integer := 0;
WRITE_WIDTH_B : integer := 0
);
port(
CASCADEOUTA  : out  std_ulogic;
CASCADEOUTB  : out  std_ulogic;
DOA          : out std_logic_vector (31 downto 0);
DOB          : out std_logic_vector (31 downto 0);
DOPA         : out std_logic_vector (3 downto 0);
DOPB         : out std_logic_vector (3 downto 0);
ADDRA        : in  std_logic_vector (14 downto 0);
ADDRB        : in  std_logic_vector (14 downto 0);
CASCADEINA   : in  std_ulogic;
CASCADEINB   : in  std_ulogic;
CLKA         : in  std_ulogic;
CLKB         : in  std_ulogic;
DIA          : in  std_logic_vector (31 downto 0);
DIB          : in  std_logic_vector (31 downto 0);
DIPA         : in  std_logic_vector (3 downto 0);
DIPB         : in  std_logic_vector (3 downto 0);
ENA          : in  std_ulogic;
ENB          : in  std_ulogic;
REGCEA       : in  std_ulogic;
REGCEB       : in  std_ulogic;
SSRA         : in  std_ulogic;
SSRB         : in  std_ulogic;
WEA          : in  std_logic_vector (3 downto 0);
WEB          : in  std_logic_vector (3 downto 0)
);
end component RAMB16;

signal odata_kvdd : std_logic_vector(31 downto 0);
signal odata_vdd25 : std_logic_vector(31 downto 0);
signal address_kvdd : std_logic_vector(14 downto 0);
signal address_vdd25 : std_logic_vector(14 downto 0);

begin

p0 : process (i_address) is
begin
	address_kvdd <= std_logic_vector(to_unsigned(to_integer(unsigned(i_address)) * 16,15));
end process p0;

p1 : process (i_address) is
begin
	address_vdd25 <= std_logic_vector(to_unsigned(((to_integer(unsigned(i_address))) * 16) + 4096,15));
end process p1;

o_data_kvdd(15 downto 0) <= odata_kvdd(15 downto 0);
o_data_vdd25(15 downto 0) <= odata_vdd25(15 downto 0);

inst_mem_kvdd : RAMB16
generic map (
DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
INIT_A => X"000000000", -- Initial values on A output port
INIT_B => X"000000000", -- Initial values on B output port
INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
READ_WIDTH_A => 18, -- Valid values are 1,2,4,9,18 or 36
READ_WIDTH_B => 18, -- Valid values are 1,2,4,9,18 or 36
SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
WRITE_MODE_A => "READ_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_MODE_B => "READ_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_WIDTH_A => 18, -- Valid values are 1,2,4,9,18 or 36
WRITE_WIDTH_B => 18, -- Valid values are 1,2,4,9,18 or 36

-- page22 11.1.1. Restoring the VDD sensor parameters
-- kvdd = (EE[0x2433] & 0xFF00) / 2^8 ; if kvdd > 127 -> kvdd = kvdd - 256 ; kvdd = kvdd * 2^5
INIT_00 => X"01e001c001a00180016001400120010000e000c000a000800060004000200000",
INIT_01 => X"03e003c003a00380036003400320030002e002c002a002800260024002200200",
INIT_02 => X"05e005c005a00580056005400520050004e004c004a004800460044004200400",
INIT_03 => X"07e007c007a00780076007400720070006e006c006a006800660064006200600",
INIT_04 => X"09e009c009a00980096009400920090008e008c008a008800860084008200800",
INIT_05 => X"0be00bc00ba00b800b600b400b200b000ae00ac00aa00a800a600a400a200a00",
INIT_06 => X"0de00dc00da00d800d600d400d200d000ce00cc00ca00c800c600c400c200c00",
INIT_07 => X"0fe00fc00fa00f800f600f400f200f000ee00ec00ea00e800e600e400e200e00",
INIT_08 => X"f1e0f1c0f1a0f180f160f140f120f100f0e0f0c0f0a0f080f060f040f020f000",
INIT_09 => X"f3e0f3c0f3a0f380f360f340f320f300f2e0f2c0f2a0f280f260f240f220f200",
INIT_0a => X"f5e0f5c0f5a0f580f560f540f520f500f4e0f4c0f4a0f480f460f440f420f400",
INIT_0b => X"f7e0f7c0f7a0f780f760f740f720f700f6e0f6c0f6a0f680f660f640f620f600",
INIT_0c => X"f9e0f9c0f9a0f980f960f940f920f900f8e0f8c0f8a0f880f860f840f820f800",
INIT_0d => X"fbe0fbc0fba0fb80fb60fb40fb20fb00fae0fac0faa0fa80fa60fa40fa20fa00",
INIT_0e => X"fde0fdc0fda0fd80fd60fd40fd20fd00fce0fcc0fca0fc80fc60fc40fc20fc00",
INIT_0f => X"ffe0ffc0ffa0ff80ff60ff40ff20ff00fee0fec0fea0fe80fe60fe40fe20fe00",
-- vdd25 = EE[0x2433] & 0x00FF ; vdd25 = (vdd25 - 256) * 2^5 - 2^13
INIT_10 => X"c1e0c1c0c1a0c180c160c140c120c100c0e0c0c0c0a0c080c060c040c020c000",
INIT_11 => X"c3e0c3c0c3a0c380c360c340c320c300c2e0c2c0c2a0c280c260c240c220c200",
INIT_12 => X"c5e0c5c0c5a0c580c560c540c520c500c4e0c4c0c4a0c480c460c440c420c400",
INIT_13 => X"c7e0c7c0c7a0c780c760c740c720c700c6e0c6c0c6a0c680c660c640c620c600",
INIT_14 => X"c9e0c9c0c9a0c980c960c940c920c900c8e0c8c0c8a0c880c860c840c820c800",
INIT_15 => X"cbe0cbc0cba0cb80cb60cb40cb20cb00cae0cac0caa0ca80ca60ca40ca20ca00",
INIT_16 => X"cde0cdc0cda0cd80cd60cd40cd20cd00cce0ccc0cca0cc80cc60cc40cc20cc00",
INIT_17 => X"cfe0cfc0cfa0cf80cf60cf40cf20cf00cee0cec0cea0ce80ce60ce40ce20ce00",
INIT_18 => X"d1e0d1c0d1a0d180d160d140d120d100d0e0d0c0d0a0d080d060d040d020d000",
INIT_19 => X"d3e0d3c0d3a0d380d360d340d320d300d2e0d2c0d2a0d280d260d240d220d200",
INIT_1a => X"d5e0d5c0d5a0d580d560d540d520d500d4e0d4c0d4a0d480d460d440d420d400",
INIT_1b => X"d7e0d7c0d7a0d780d760d740d720d700d6e0d6c0d6a0d680d660d640d620d600",
INIT_1c => X"d9e0d9c0d9a0d980d960d940d920d900d8e0d8c0d8a0d880d860d840d820d800",
INIT_1d => X"dbe0dbc0dba0db80db60db40db20db00dae0dac0daa0da80da60da40da20da00",
INIT_1e => X"dde0ddc0dda0dd80dd60dd40dd20dd00dce0dcc0dca0dc80dc60dc40dc20dc00",
INIT_1f => X"dfe0dfc0dfa0df80df60df40df20df00dee0dec0dea0de80de60de40de20de00",

INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
)
port map (
CASCADEOUTA => open, -- 1-bit cascade output
CASCADEOUTB => open, -- 1-bit cascade output
DOA => odata_kvdd, -- 32-bit A port Data Output
DOB => odata_vdd25, -- 32-bit B port Data Output
DOPA => open, -- 4-bit A port Parity Output
DOPB => open, -- 4-bit B port Parity Output
ADDRA => address_kvdd, -- 15-bit A port Address Input
ADDRB => address_vdd25, -- 15-bit B port Address Input
CASCADEINA => '0', -- 1-bit cascade A input
CASCADEINB => '0', -- 1-bit cascade B input
CLKA => i_clock, -- Port A Clock
CLKB => i_clock, -- Port B Clock
DIA => (others => '0'), -- 32-bit A port Data Input
DIB => (others => '0'), -- 32-bit B port Data Input
DIPA => (others => '0'), -- 4-bit A port parity Input
DIPB => (others => '0'), -- 4-bit B port parity Input
ENA => '1', -- 1-bit A port Enable Input
ENB => '1', -- 1-bit B port Enable Input
REGCEA => '1', -- 1-bit A port register enable input
REGCEB => '1', -- 1-bit B port register enable input
SSRA => i_reset, -- 1-bit A port Synchronous Set/Reset Input
SSRB => i_reset, -- 1-bit B port Synchronous Set/Reset Input
WEA => (others => '0'), -- 4-bit A port Write Enable Input
WEB => (others => '0') -- 4-bit B port Write Enable Input
);

--RAMB16
--generic map (
--DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
--DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
--INIT_A => X"000000000", -- Initial values on A output port
--INIT_B => X"000000000", -- Initial values on B output port
--INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
--INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
--RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--READ_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36
--READ_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
--SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
--SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
--WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
--WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
--WRITE_WIDTH_A => 2, -- Valid values are 1,2,4,9,18 or 36
--WRITE_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
--INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
--INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
--)
--port map (
--CASCADEOUTA => CASCADEOUTA, -- 1-bit cascade output
--CASCADEOUTB => CASCADEOUTB, -- 1-bit cascade output
--DOA => DOA, -- 32-bit A port Data Output
--DOB => DOB, -- 32-bit B port Data Output
--DOPA => DOPA, -- 4-bit A port Parity Output
--DOPB => DOPB, -- 4-bit B port Parity Output
--ADDRA => ADDRA, -- 15-bit A port Address Input
--ADDRB => ADDRB, -- 15-bit B port Address Input
--CASCADEINA => CASCADEINA, -- 1-bit cascade A input
--CASCADEINB => CASCADEINB, -- 1-bit cascade B input
--CLKA => CLKA, -- Port A Clock
--CLKB => CLKB, -- Port B Clock
--DIA => DIA, -- 32-bit A port Data Input
--DIB => DIB, -- 32-bit B port Data Input
--DIPA => DIPA, -- 4-bit A port parity Input
--DIPB => DIPB, -- 4-bit B port parity Input
--ENA => ENA, -- 1-bit A port Enable Input
--ENB => ENB, -- 1-bit B port Enable Input
--REGCEA => REGCEA, -- 1-bit A port register enable input
--REGCEB => REGCEB, -- 1-bit B port register enable input
--SSRA => SSRA, -- 1-bit A port Synchronous Set/Reset Input
--SSRB => SSRB, -- 1-bit B port Synchronous Set/Reset Input
--WEA => WEA, -- 4-bit A port Write Enable Input
--WEB => WEB -- 4-bit B port Write Enable Input
--);

end Behavioral;
