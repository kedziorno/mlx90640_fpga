----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:51:51 12/19/2022 
-- Design Name: 
-- Module Name:    mem_16bit_address - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mem_ramb16_16bit_address is
port (
O_CASCADEOUTA  : out std_ulogic;
O_CASCADEOUTB  : out std_ulogic;
O_DOA          : out std_logic_vector (31 downto 0);
O_DOB          : out std_logic_vector (31 downto 0);
O_DOPA         : out std_logic_vector (3 downto 0);
O_DOPB         : out std_logic_vector (3 downto 0);
I_ADDRA        : in  std_logic_vector (15 downto 0); -- 16bit
I_ADDRB        : in  std_logic_vector (15 downto 0); -- 16bit
I_CASCADEINA   : in  std_ulogic;
I_CASCADEINB   : in  std_ulogic;
I_CLKA         : in  std_ulogic;
I_CLKB         : in  std_ulogic;
I_DIA          : in  std_logic_vector (31 downto 0);
I_DIB          : in  std_logic_vector (31 downto 0);
I_DIPA         : in  std_logic_vector (3 downto 0);
I_DIPB         : in  std_logic_vector (3 downto 0);
I_ENA          : in  std_ulogic;
I_ENB          : in  std_ulogic;
I_REGCEA       : in  std_ulogic;
I_REGCEB       : in  std_ulogic;
I_SSRA         : in  std_ulogic;
I_SSRB         : in  std_ulogic;
I_WEA          : in  std_logic_vector (3 downto 0);
I_WEB          : in  std_logic_vector (3 downto 0)
end entity mem_ramb16_16bit_address;

architecture Behavioral of mem_16bit_address is

component RAMB16 is
generic (
DOA_REG : integer := 0 ;
DOB_REG : integer := 0 ;
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_A : bit_vector := X"000000000";
INIT_B : bit_vector := X"000000000";
INIT_FILE : string := "NONE";
INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INVERT_CLK_DOA_REG : boolean := false;
INVERT_CLK_DOB_REG : boolean := false;
RAM_EXTENSION_A : string := "NONE";
RAM_EXTENSION_B : string := "NONE";
READ_WIDTH_A : integer := 0;
READ_WIDTH_B : integer := 0;
SIM_COLLISION_CHECK : string := "ALL";
SRVAL_A  : bit_vector := X"000000000";
SRVAL_B  : bit_vector := X"000000000";
WRITE_MODE_A : string := "WRITE_FIRST";
WRITE_MODE_B : string := "WRITE_FIRST";
WRITE_WIDTH_A : integer := 0;
WRITE_WIDTH_B : integer := 0
);
port(
CASCADEOUTA  : out  std_ulogic;
CASCADEOUTB  : out  std_ulogic;
DOA          : out std_logic_vector (31 downto 0);
DOB          : out std_logic_vector (31 downto 0);
DOPA         : out std_logic_vector (3 downto 0);
DOPB         : out std_logic_vector (3 downto 0);
ADDRA        : in  std_logic_vector (14 downto 0);
ADDRB        : in  std_logic_vector (14 downto 0);
CASCADEINA   : in  std_ulogic;
CASCADEINB   : in  std_ulogic;
CLKA         : in  std_ulogic;
CLKB         : in  std_ulogic;
DIA          : in  std_logic_vector (31 downto 0);
DIB          : in  std_logic_vector (31 downto 0);
DIPA         : in  std_logic_vector (3 downto 0);
DIPB         : in  std_logic_vector (3 downto 0);
ENA          : in  std_ulogic;
ENB          : in  std_ulogic;
REGCEA       : in  std_ulogic;
REGCEB       : in  std_ulogic;
SSRA         : in  std_ulogic;
SSRB         : in  std_ulogic;
WEA          : in  std_logic_vector (3 downto 0);
WEB          : in  std_logic_vector (3 downto 0)
);
end component RAMB16;

signal mux : std_logic;

signal CASCADEOUTA_lo,CASCADEOUTB_lo,CASCADEINA_lo,CASCADEINB_lo,CLKA_lo,CLKB_lo,ENA_lo,ENB_lo,REGCEA_lo,REGCEB_lo,SSRA_lo,SSRB_lo : std_logic;
signal DOA_lo,DOB_lo,DIA_lo,DIB_lo : std_logic_vector(31 downto 0);
signal DOPA_lo,DOPB_lo,DIPA_lo,DIPB_lo,WEA_lo,WEB_lo : std_logic_vector(3 downto 0);
signal ADDRA_lo,ADDRB_lo : std_logic_vector(14 downto 0);

signal CASCADEOUTA_hi,CASCADEOUTB_hi,CASCADEINA_hi,CASCADEINB_hi,CLKA_hi,CLKB_hi,ENA_hi,ENB_hi,REGCEA_hi,REGCEB_hi,SSRA_hi,SSRB_hi : std_logic;
signal DOA_hi,DOB_hi,DIA_hi,DIB_hi : std_logic_vector(31 downto 0);
signal DOPA_hi,DOPB_hi,DIPA_hi,DIPB_hi,WEA_hi,WEB_hi : std_logic_vector(3 downto 0);
signal ADDRA_hi,ADDRB_hi : std_logic_vector(14 downto 0);

begin

mux <= '1' when (I_ADDRA(15) = '1' or I_ADDRB(15) = '1') else '0';

O_CASCADEOUTA <= CASCADEOUTA_lo when mux = '0' else CASCADEOUTA_hi when mux = '1' else '0';
O_CASCADEOUTB <= CASCADEOUTB_lo when mux = '0' else CASCADEOUTB_hi when mux = '1' else '0';
O_DOA <= DOA_lo when mux = '0' else DOA_hi when mux = '1' else (others => '0');
O_DOB <= DOB_lo when mux = '0' else DOB_hi when mux = '1' else (others => '0');
O_DOPA <= DOPA_lo when mux = '0' else DOPA_hi when mux = '1' else (others => '0');
O_DOPB <= DOPB_lo when mux = '0' else DOPB_hi when mux = '1' else (others => '0');
ADDRA_lo <= I_ADDRA when mux = '0' else (others => '0');
ADDRA_hi <= I_ADDRA when mux = '1' else (others => '0');
ADDRB_lo <= I_ADDRB when mux = '0' else (others => '0');
ADDRB_hi <= I_ADDRB when mux = '1' else (others => '0');
CASCADEINA_lo <= I_CASCADEINA when mux = '0' else '0';
CASCADEINA_hi <= I_CASCADEINA when mux = '1' else '0';
CASCADEINB_lo <= I_CASCADEINB when mux = '0' else '0';
CASCADEINB_hi <= I_CASCADEINB when mux = '1' else '0';
CLKA_lo <= I_CLKA when mux = '0' else '0';
CLKA_hi <= I_CLKA when mux = '1' else '0';
CLKB_lo <= I_CLKB when mux = '0' else '0';
CLKB_hi <= I_CLKB when mux = '1' else '0';
DIA_lo <= I_DIA when mux = '0' else (others => '0');
DIA_hi <= I_DIA when mux = '1' else (others => '0');
DIB_lo <= I_DIB when mux = '0' else (others => '0');
DIB_hi <= I_DIB when mux = '1' else (others => '0');
DIPA_lo <= I_DIPA when mux = '0' else (others => '0');
DIPA_hi <= I_DIPA when mux = '1' else (others => '0');
DIPB_lo <= I_DIPB when mux = '0' else (others => '0');
DIPB_hi <= I_DIPB when mux = '1' else (others => '0');
ENA_lo <= I_ENA when mux = '0' else '0';
ENA_hi <= I_ENA when mux = '1' else '0';
ENB_lo <= I_ENB when mux = '0' else '0';
ENB_hi <= I_ENB when mux = '1' else '0';
REGCEA_lo <= I_REGCEA when mux = '0' else '0';
REGCEA_hi <= I_REGCEA when mux = '1' else '0';
REGCEB_lo <= I_REGCEB when mux = '0' else '0';
REGCEB_hi <= I_REGCEB when mux = '1' else '0';
SSRA_lo <= I_SSRA when mux = '0' else '0';
SSRA_hi <= I_SSRA when mux = '1' else '0';
SSRB_lo <= I_SSRB when mux = '0' else '0';
SSRB_hi <= I_SSRB when mux = '1' else '0';
WEA_lo <= I_WEA when mux = '0' else (others => '0');
WEA_hi <= I_WEA when mux = '1' else (others => '0');
WEB_lo <= I_WEB when mux = '0' else (others => '0');
WEB_hi <= I_WEB when mux = '1' else (others => '0');

inst_ramb16_hi : RAMB16
generic map (
DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
INIT_A => X"000000000", -- Initial values on A output port
INIT_B => X"000000000", -- Initial values on B output port
INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
READ_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36
READ_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_WIDTH_A => 2, -- Valid values are 1,2,4,9,18 or 36
WRITE_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
)
port map (
CASCADEOUTA => CASCADEOUTA_hi, -- 1-bit cascade output
CASCADEOUTB => CASCADEOUTB_hi, -- 1-bit cascade output
DOA => DOA_hi, -- 32-bit A port Data Output
DOB => DOB_hi, -- 32-bit B port Data Output
DOPA => DOPA_hi, -- 4-bit A port Parity Output
DOPB => DOPB_hi, -- 4-bit B port Parity Output
ADDRA => ADDRA_hi, -- 15-bit A port Address Input
ADDRB => ADDRB_hi, -- 15-bit B port Address Input
CASCADEINA => CASCADEINA_hi, -- 1-bit cascade A input
CASCADEINB => CASCADEINB_hi, -- 1-bit cascade B input
CLKA => CLKA_hi, -- Port A Clock
CLKB => CLKB_hi, -- Port B Clock
DIA => DIA_hi, -- 32-bit A port Data Input
DIB => DIB_hi, -- 32-bit B port Data Input
DIPA => DIPA_hi, -- 4-bit A port parity Input
DIPB => DIPB_hi, -- 4-bit B port parity Input
ENA => ENA_hi, -- 1-bit A port Enable Input
ENB => ENB_hi, -- 1-bit B port Enable Input
REGCEA => REGCEA_hi, -- 1-bit A port register enable input
REGCEB => REGCEB_hi, -- 1-bit B port register enable input
SSRA => SSRA_hi, -- 1-bit A port Synchronous Set/Reset Input
SSRB => SSRB_hi, -- 1-bit B port Synchronous Set/Reset Input
WEA => WEA_hi, -- 4-bit A port Write Enable Input
WEB => WEB_hi -- 4-bit B port Write Enable Input
);

inst_ramb16_lo : RAMB16
generic map (
DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
INIT_A => X"000000000", -- Initial values on A output port
INIT_B => X"000000000", -- Initial values on B output port
INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
READ_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36
READ_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
SRVAL_A => X"000000000", -- Port A ouput value upon SSR assertion
SRVAL_B => X"000000000", -- Port B ouput value upon SSR assertion
WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
WRITE_WIDTH_A => 2, -- Valid values are 1,2,4,9,18 or 36
WRITE_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
)
port map (
CASCADEOUTA => CASCADEOUTA_lo, -- 1-bit cascade output
CASCADEOUTB => CASCADEOUTB_lo, -- 1-bit cascade output
DOA => DOA_lo, -- 32-bit A port Data Output
DOB => DOB_lo, -- 32-bit B port Data Output
DOPA => DOPA_lo, -- 4-bit A port Parity Output
DOPB => DOPB_lo, -- 4-bit B port Parity Output
ADDRA => ADDRA_lo, -- 15-bit A port Address Input
ADDRB => ADDRB_lo, -- 15-bit B port Address Input
CASCADEINA => CASCADEINA_lo, -- 1-bit cascade A input
CASCADEINB => CASCADEINB_lo, -- 1-bit cascade B input
CLKA => CLKA_lo, -- Port A Clock
CLKB => CLKB_lo, -- Port B Clock
DIA => DIA_lo, -- 32-bit A port Data Input
DIB => DIB_lo, -- 32-bit B port Data Input
DIPA => DIPA_lo, -- 4-bit A port parity Input
DIPB => DIPB_lo, -- 4-bit B port parity Input
ENA => ENA_lo, -- 1-bit A port Enable Input
ENB => ENB_lo, -- 1-bit B port Enable Input
REGCEA => REGCEA_lo, -- 1-bit A port register enable input
REGCEB => REGCEB_lo, -- 1-bit B port register enable input
SSRA => SSRA_lo, -- 1-bit A port Synchronous Set/Reset Input
SSRB => SSRB_lo, -- 1-bit B port Synchronous Set/Reset Input
WEA => WEA_lo, -- 4-bit A port Write Enable Input
WEB => WEB_lo -- 4-bit B port Write Enable Input
);

end Behavioral;
