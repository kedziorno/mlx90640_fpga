----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:39:33 08/24/2024 
-- Design Name: 
-- Module Name:    tfm_mock - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tfm_mock is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_run : in std_logic;

i2c_mem_ena : out STD_LOGIC;
i2c_mem_addra : out STD_LOGIC_VECTOR(11 DOWNTO 0);
i2c_mem_douta : in STD_LOGIC_VECTOR(7 DOWNTO 0);

o_rdy : out std_logic;

i_addr : in std_logic_vector(9 downto 0);
o_do : out std_logic_vector(31 downto 0)
);
end tfm_mock;

architecture Behavioral of tfm_mock is

COMPONENT mem_ramb16_s36_x2
generic (
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0a : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0b : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0c : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0d : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0e : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0f : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
);
PORT(
DO : OUT  std_logic_vector(31 downto 0);
DOP : OUT  std_logic_vector(3 downto 0);
ADDR : IN  std_logic_vector(9 downto 0);
CLK : IN  std_logic;
DI : IN  std_logic_vector(31 downto 0);
DIP : IN  std_logic_vector(3 downto 0);
EN : IN  std_logic;
SSR : IN  std_logic;
WE : IN  std_logic
);
END COMPONENT mem_ramb16_s36_x2;

begin

p0 : process (i_clock, i_reset) is
type states is (a, b);
variable state : states;
begin
  if (i_reset = '1') then
    o_rdy <= '0';
    state := a;
  elsif (rising_edge (i_clock)) then
    case (state) is
      when a =>
        o_rdy <= '0';
        if (i_run = '1') then
          state := b;
        else
          state := a;
        end if;
      when b =>
        o_rdy <= '1';
        state := b;
    end case;
  end if;
end process p0;

i2c_mem_ena <= '0';
i2c_mem_addra <= (others => '0');

inst_calculated_to : mem_ramb16_s36_x2 
GENERIC MAP (
INIT_00 => X"41E2EB5041E57D4041E3B2D041E2EB5041E23AF041E1CB2041DE70907FC00000",
INIT_01 => X"41DFE25041E5F64041E27FE041E3300041E04D1041E52DA041E1E15041E2D6B0",
INIT_02 => X"41E1771041E5756041E64DB041E976D041E2006041E5120041E4652041E28430",
INIT_03 => X"41E9464041ED93D041E8A15041E7437041E41E9041E7746041E5D07041E8F7A0",
INIT_04 => X"41E08A7041E35DB041E4C7B041E488F041E1B6A041E2DE1041E5867041E7BA90",
INIT_05 => X"41E2C70041DF1DE041E1F04041E63A4041E0049041E16CC041E16CC041E2C280",
INIT_06 => X"41E6736041E5257041E753E041E315E041E4E21041E4DC9041E2444041E129A0",
INIT_07 => X"41E85D3041E857B041E54BA041E73E3041E4FC2041E50B6041E713F041E51670",
INIT_08 => X"41E09AC041E04DA041E6541041E4198041E1749041E483E041E50B4041E4B530",
INIT_09 => X"41E393E041E1C77041E4F61041E3790041E1D01041E3D6D041E3D02041E2BA90",
INIT_0a => X"41E3799041E445C041E37EB041E89B8041E0CD7041E34FA041E243C041E51C70",
INIT_0b => X"41E3051041E5A73041E59E5041E8DA6041E2D23041E6DCA041E473A041E68650",
INIT_0c => X"41E4D72041E29CB041E214A041E3A72041E28E6041E3A74041E18E9041E41260",
INIT_0d => X"41E4717041E2FC6041E2AEC041E2D81041E11F5041E3732041E3223041E1A720",
INIT_0e => X"41E47D6041E573F041E7550041E4FC0041E3BA1041E2A64041E2AE0041E2FA80",
INIT_0f => X"41E89B5041E297F041E4B9F041E6908041E4019041E434F041E73B0041E5FD10",
INIT_10 => X"41E2409041E43EA041E4B18041E2DEA041E2E6E041E66D5041E2EE8041E1F630",
INIT_11 => X"41DFA22041E697F041E2337041E4492041E3382041E2599041E612D041E59BE0",
INIT_12 => X"41E4234041E53D0041E7619041E2CAB041E420D041E2D0E041E2703041E3AEC0",
INIT_13 => X"41DCAB9041E7E53041E6BBD041E6934041E38C1041E85AC041E3AA2041E57890",
INIT_14 => X"41E30B0041E7EFA041E39C9041E3EF6041E055F041E3FE9041E1895041E139D0",
INIT_15 => X"41E325C041E1478041E2FA9041E37B2041E5994041E69F9041E3654041ECCF80",
INIT_16 => X"41E4EEE041E4807041E677C041D107A041E661A041E3C09041E2AEC041E6A020",
INIT_17 => X"41E2038041E2718041E50D0041E62BA041E6114041E58AF041E4945041E4B8C0",
INIT_18 => X"41E69DB041E4B8A041E4BC9041E598B041E3C31041E3115041E2ECE041E48EB0",
INIT_19 => X"41E3A15041E3585041E6F0C041E6DDA041EED60041EBA62041F8D71041EA34A0",
INIT_1a => X"41E359E041E8555041E20F0041E5CA3041E1572041E5E3E041E272E041E58730",
INIT_1b => X"41DA1AE041E769B041E29E3041E445D041E4E15041E37DF041E4D62041E09A70",
INIT_1c => X"41E2B2C041E5D29041E0E5F041E5441041E2A3F041E53E0041E38E3041E421B0",
INIT_1d => X"41E5DD0041E5AAD041E60ED041EEA32041F0F1D041FAED7041ED40B041FD3B70",
INIT_1e => X"41E20A0041E4124041E4421041E3CC6041E3357041E3AD4041E3411041E50B90",
INIT_1f => X"41DFC6E041E02F0041E6F07041E624E041E41DC041E44A8041E3E0A041E4D800",
INIT_20 => X"41F2906041E73E3041E8292041E33B3041E4530041E57D7041E3E32041E16610",
INIT_21 => X"41EB8D1041EB42A041FA4AE041FB4AB0420069F04201C170420265F041F4F190",
INIT_22 => X"41E4A2D041E62BB041E1C13041E5EB2041E3E46041E4E6B041E4EE1041E1D110",
INIT_23 => X"41D9974041E6829041E30B8041E50BC041E27CB041E6678041E2CDA041E4A250",
INIT_24 => X"41E86AF041F46CA041E44A4041E7C7C041E0565041E31A7041E2D95041E47FD0",
INIT_25 => X"41EF325041F77CD041FAEA404202F0684200ABA04202C1E041FF9E9042038F78",
INIT_26 => X"41E575A041E3C4F041E7269041E597F041E3268041E551D041E5769041E9FE50",
INIT_27 => X"41E3334041DD4E5041E3EC6041E64AF041E54AE041E21C2041E3910041E2AD90",
INIT_28 => X"4202457841ECE9F041EC080041E686D041E6F2D041E60D8041E641B041E570B0",
INIT_29 => X"4200C9684200A1B04202AFB04202A9184203FF804203CDF042063E304201A4E8",
INIT_2a => X"41E248E041E3B89041E5297041E3903041E4B29041EAD0B041F336C041F34900",
INIT_2b => X"41E17E5041E534F041E42E2041E5D81041E3E07041E6E7C041E3DFF041E579A0",
INIT_2c => X"41F3F1204201365041E6B5B041EC6B0041E4862041E1F92041E349B041E6E180",
INIT_2d => X"42002A304200E3484203AAC84203A1584204F7C04206579842052AA842093078",
INIT_2e => X"41E5C3F041DFA9F041E463E041E2D5C041E969A041ED0E2041F6A3A041FF0C80",
INIT_2f => X"41E469F041E5A6D041E4632041E5013041E642F041E404C041E4252041E1A9F0",
INIT_30 => X"420618D041F7603041F8DB6041E8436041E39C7041E2593041E2CBD041E44010",
INIT_31 => X"420186004202C9184202AFB0420619C042076CE84208E188420A3E904206C8A8",
INIT_32 => X"41E4011041E5066041E5C7C041E84E4041E79B0041FA1C2041FD5540420131F0",
INIT_33 => X"41E348B041E5C1C041E1F2D041E48BC041E3705041E366B041E2E9C041E396A0",
INIT_34 => X"42014FB04202B23041EA29F041F632F041E28ED041E6A18041E3FD0041E74FB0",
INIT_35 => X"420249F0420321B84205B9884205D8C04209C8284207C9B8420874384207BD90",
INIT_36 => X"41E1ADE041E4006041E650E041E621D041F50CB041EB14C0420268B841FDB8F0",
INIT_37 => X"41E4206041E4AA4041E5DFA041E6F40041E419E041E26C3041E45D9041E46250",
INIT_38 => X"42026FC04202586841FFEE4041EC2B7041E6E90041E59E5041E66EB041E3ED30",
INIT_39 => X"4202E478420578104202DBC842061EF04204D1604209A49842055EF84206CC80",
INIT_3a => X"41E2030041E6BB3041E5808041E7F58041E73B7041F5551041F6478042021388",
INIT_3b => X"41E312D041E71A7041E422E041E604C041E437D041E513A041E4998041E46270",
INIT_3c => X"420361004202B92841F1B20041FCBC0041E810D041E83E3041E3A52041E37060",
INIT_3d => X"4202FF1042025670420466484203D31842070EA84202FDD04205B4884202FCD8",
INIT_3e => X"41E2171041E6030041E72CC041E439D041EAD52041E7575042024CB841FAFBE0",
INIT_3f => X"41E73B3041E5BE4041E4134041E6E52041E3111041E6E8E041E2E42041E38C60",
INIT_40 => X"420255B84204AFE841FB288041F79C0041EC08E041ED2C8041EDDFB041E99860",
INIT_41 => X"42016768420653284205AEE8420587904204BB00420711A84204E9D042057EC8",
INIT_42 => X"41E7F9A041ED55F041E8B91041EA99B041E9178041F1CA6041F15C404204CCC8",
INIT_43 => X"41F0EE6041EF975041EFCD0041F1866041F21EA041EC0F0041E9D92041E851C0",
INIT_44 => X"42013C5041F7D7C041F41E1041EC3BA041E88C8041E5DA2041E2A9D041E1BE30",
INIT_45 => X"4202FAF041FED2C04203AC38420274F842018368420195D04201425841FEED40",
INIT_46 => X"41E43B6041E1772041E36C9041E5A22041E5A45041E3C97041F91B0041F0FD00",
INIT_47 => X"41E8174041E6683041EE368041F2B3B041E6232041EBA9F041E5F06041E4C4E0",
INIT_48 => X"41EB899041EF415041E62F8041E9ED5041E35F6041E52EB041E4A5B041E3FC60",
INIT_49 => X"41F114E04202A4D8420149D04201581841FF5F904201CB6041F67A2041FDF1F0",
INIT_4a => X"41E2B1C041E4C07041E563D041E568A041E42CC041EA6D8041E7506041FA0890",
INIT_4b => X"41EEA83041FCC9504201595041FA12B041FA448041EA676041E62EA041E851C0",
INIT_4c => X"41EE392041E6929041E511C041E412D041E44AF041E27FA041E1A52041E74D00",
INIT_4d => X"4200483041F484D042003A3841FDA4B041FD5E1041F3EBA041F443B041EB5F50",
INIT_4e => X"41E6289041E3064041E267F041E49F3041E46FF041E1FAA041EDA01041E7A270",
INIT_4f => X"4200D2284201F1F042025AF842034E7841EF234041F7106041E6321041E8B070",
INIT_50 => X"41E57E8041E3A23041E3552041E5E5F041E3BF0041E2B0C041E4275041E44620",
INIT_51 => X"41EA367041FA89A041F1C7D041F8980041ECF31041EF027041E663A041EA71B0",
INIT_52 => X"41E3A24041E43D7041E5024041E4ED4041E4770041E4C1D041E1840041ED4300",
INIT_53 => X"42001B08420913D0420808984201DCE042015A3841F5523041EE498041E5C6E0",
INIT_54 => X"41E4BBB041E3D30041E20B3041E51E5041E12DE041E35FF041E310C041E798D0",
INIT_55 => X"41F2A14041E752D041F3B78041E8AC7041E8A69041E7F40041E55A3041E6FB10",
INIT_56 => X"41E293D041E2F22041E5173041E5A8E041E2FB9041E217E041E695F041E6AA20",
INIT_57 => X"4204F3A84202D5D8420522B04207679841FB0C7041FD813041E5441041EF7D00",
INIT_58 => X"41E2325041E754B041E3EBB041E44C0041E0734041E30DE041E2181041E49400",
INIT_59 => X"41E3FA9041E8736041E4CA6041E780B041E3B2B041E4549041E359D041E5BFB0",
INIT_5a => X"41E6D74041E7482041E3337041E2E64041E3206041E7478041E4351041E8F640",
INIT_5b => X"41F2727042040C184204F0C0420489D84202093041FFEEA041FA2CA041E902E0",
INIT_5c => X"41E2E84041E339E041E33E3041E38C8041E27DC041E2B24041E1A86041E24AF0",
INIT_5d => X"41E7ED5041E3531041E575B041E4284041E2D59041E599D041E1573041E26D60",
INIT_5e => X"41E3C43041E49A4041E3A45041E4539041E1F68041DFFAB041E4A1F041E522F0",
INIT_5f => X"42001DA841F8CEF04202320842045B1842028E00420280C041F1B11041FD3C00"
)
PORT MAP (
DO => o_do,
DOP => open,
ADDR => i_addr,
CLK => i_clock,
DI => (others => '0'),
DIP => (others => '0'),
EN => '1',
SSR => i_reset,
WE => '0'
);

end Behavioral;

