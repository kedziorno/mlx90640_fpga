----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:39:33 08/24/2024 
-- Design Name: 
-- Module Name:    tfm_mock - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tfm_mock is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_run : in std_logic;

i2c_mem_ena : out STD_LOGIC;
i2c_mem_addra : out STD_LOGIC_VECTOR(11 DOWNTO 0);
i2c_mem_douta : in STD_LOGIC_VECTOR(7 DOWNTO 0);

o_rdy : out std_logic;

i_addr : in std_logic_vector(9 downto 0);
o_do : out std_logic_vector(31 downto 0)
);
end tfm_mock;

architecture Behavioral of tfm_mock is

COMPONENT mem_ramb16_s36_x2
generic (
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0a : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0b : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0c : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0d : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0e : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0f : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
);
PORT(
DO : OUT  std_logic_vector(31 downto 0);
DOP : OUT  std_logic_vector(3 downto 0);
ADDR : IN  std_logic_vector(9 downto 0);
CLK : IN  std_logic;
DI : IN  std_logic_vector(31 downto 0);
DIP : IN  std_logic_vector(3 downto 0);
EN : IN  std_logic;
SSR : IN  std_logic;
WE : IN  std_logic
);
END COMPONENT mem_ramb16_s36_x2;

begin

p0 : process (i_clock, i_reset) is
type states is (a, b);
variable state : states;
begin
  if (i_reset = '1') then
    o_rdy <= '0';
    state := a;
  elsif (rising_edge (i_clock)) then
    case (state) is
      when a =>
        o_rdy <= '0';
        if (i_run = '1') then
          state := b;
        else
          state := a;
        end if;
      when b =>
        o_rdy <= '1';
        state := b;
    end case;
  end if;
end process p0;

i2c_mem_ena <= '0';
i2c_mem_addra <= (others => '0');

inst_calculated_to : mem_ramb16_s36_x2
--GENERIC MAP ( -- XXX temperatures
--INIT_00 => X"41E2EB5041E57D4041E3B2D041E2EB5041E23AF041E1CB2041DE70907FC00000",
--INIT_01 => X"41DFE25041E5F64041E27FE041E3300041E04D1041E52DA041E1E15041E2D6B0",
--INIT_02 => X"41E1771041E5756041E64DB041E976D041E2006041E5120041E4652041E28430",
--INIT_03 => X"41E9464041ED93D041E8A15041E7437041E41E9041E7746041E5D07041E8F7A0",
--INIT_04 => X"41E08A7041E35DB041E4C7B041E488F041E1B6A041E2DE1041E5867041E7BA90",
--INIT_05 => X"41E2C70041DF1DE041E1F04041E63A4041E0049041E16CC041E16CC041E2C280",
--INIT_06 => X"41E6736041E5257041E753E041E315E041E4E21041E4DC9041E2444041E129A0",
--INIT_07 => X"41E85D3041E857B041E54BA041E73E3041E4FC2041E50B6041E713F041E51670",
--INIT_08 => X"41E09AC041E04DA041E6541041E4198041E1749041E483E041E50B4041E4B530",
--INIT_09 => X"41E393E041E1C77041E4F61041E3790041E1D01041E3D6D041E3D02041E2BA90",
--INIT_0a => X"41E3799041E445C041E37EB041E89B8041E0CD7041E34FA041E243C041E51C70",
--INIT_0b => X"41E3051041E5A73041E59E5041E8DA6041E2D23041E6DCA041E473A041E68650",
--INIT_0c => X"41E4D72041E29CB041E214A041E3A72041E28E6041E3A74041E18E9041E41260",
--INIT_0d => X"41E4717041E2FC6041E2AEC041E2D81041E11F5041E3732041E3223041E1A720",
--INIT_0e => X"41E47D6041E573F041E7550041E4FC0041E3BA1041E2A64041E2AE0041E2FA80",
--INIT_0f => X"41E89B5041E297F041E4B9F041E6908041E4019041E434F041E73B0041E5FD10",
--INIT_10 => X"41E2409041E43EA041E4B18041E2DEA041E2E6E041E66D5041E2EE8041E1F630",
--INIT_11 => X"41DFA22041E697F041E2337041E4492041E3382041E2599041E612D041E59BE0",
--INIT_12 => X"41E4234041E53D0041E7619041E2CAB041E420D041E2D0E041E2703041E3AEC0",
--INIT_13 => X"41DCAB9041E7E53041E6BBD041E6934041E38C1041E85AC041E3AA2041E57890",
--INIT_14 => X"41E30B0041E7EFA041E39C9041E3EF6041E055F041E3FE9041E1895041E139D0",
--INIT_15 => X"41E325C041E1478041E2FA9041E37B2041E5994041E69F9041E3654041ECCF80",
--INIT_16 => X"41E4EEE041E4807041E677C041D107A041E661A041E3C09041E2AEC041E6A020",
--INIT_17 => X"41E2038041E2718041E50D0041E62BA041E6114041E58AF041E4945041E4B8C0",
--INIT_18 => X"41E69DB041E4B8A041E4BC9041E598B041E3C31041E3115041E2ECE041E48EB0",
--INIT_19 => X"41E3A15041E3585041E6F0C041E6DDA041EED60041EBA62041F8D71041EA34A0",
--INIT_1a => X"41E359E041E8555041E20F0041E5CA3041E1572041E5E3E041E272E041E58730",
--INIT_1b => X"41DA1AE041E769B041E29E3041E445D041E4E15041E37DF041E4D62041E09A70",
--INIT_1c => X"41E2B2C041E5D29041E0E5F041E5441041E2A3F041E53E0041E38E3041E421B0",
--INIT_1d => X"41E5DD0041E5AAD041E60ED041EEA32041F0F1D041FAED7041ED40B041FD3B70",
--INIT_1e => X"41E20A0041E4124041E4421041E3CC6041E3357041E3AD4041E3411041E50B90",
--INIT_1f => X"41DFC6E041E02F0041E6F07041E624E041E41DC041E44A8041E3E0A041E4D800",
--INIT_20 => X"41F2906041E73E3041E8292041E33B3041E4530041E57D7041E3E32041E16610",
--INIT_21 => X"41EB8D1041EB42A041FA4AE041FB4AB0420069F04201C170420265F041F4F190",
--INIT_22 => X"41E4A2D041E62BB041E1C13041E5EB2041E3E46041E4E6B041E4EE1041E1D110",
--INIT_23 => X"41D9974041E6829041E30B8041E50BC041E27CB041E6678041E2CDA041E4A250",
--INIT_24 => X"41E86AF041F46CA041E44A4041E7C7C041E0565041E31A7041E2D95041E47FD0",
--INIT_25 => X"41EF325041F77CD041FAEA404202F0684200ABA04202C1E041FF9E9042038F78",
--INIT_26 => X"41E575A041E3C4F041E7269041E597F041E3268041E551D041E5769041E9FE50",
--INIT_27 => X"41E3334041DD4E5041E3EC6041E64AF041E54AE041E21C2041E3910041E2AD90",
--INIT_28 => X"4202457841ECE9F041EC080041E686D041E6F2D041E60D8041E641B041E570B0",
--INIT_29 => X"4200C9684200A1B04202AFB04202A9184203FF804203CDF042063E304201A4E8",
--INIT_2a => X"41E248E041E3B89041E5297041E3903041E4B29041EAD0B041F336C041F34900",
--INIT_2b => X"41E17E5041E534F041E42E2041E5D81041E3E07041E6E7C041E3DFF041E579A0",
--INIT_2c => X"41F3F1204201365041E6B5B041EC6B0041E4862041E1F92041E349B041E6E180",
--INIT_2d => X"42002A304200E3484203AAC84203A1584204F7C04206579842052AA842093078",
--INIT_2e => X"41E5C3F041DFA9F041E463E041E2D5C041E969A041ED0E2041F6A3A041FF0C80",
--INIT_2f => X"41E469F041E5A6D041E4632041E5013041E642F041E404C041E4252041E1A9F0",
--INIT_30 => X"420618D041F7603041F8DB6041E8436041E39C7041E2593041E2CBD041E44010",
--INIT_31 => X"420186004202C9184202AFB0420619C042076CE84208E188420A3E904206C8A8",
--INIT_32 => X"41E4011041E5066041E5C7C041E84E4041E79B0041FA1C2041FD5540420131F0",
--INIT_33 => X"41E348B041E5C1C041E1F2D041E48BC041E3705041E366B041E2E9C041E396A0",
--INIT_34 => X"42014FB04202B23041EA29F041F632F041E28ED041E6A18041E3FD0041E74FB0",
--INIT_35 => X"420249F0420321B84205B9884205D8C04209C8284207C9B8420874384207BD90",
--INIT_36 => X"41E1ADE041E4006041E650E041E621D041F50CB041EB14C0420268B841FDB8F0",
--INIT_37 => X"41E4206041E4AA4041E5DFA041E6F40041E419E041E26C3041E45D9041E46250",
--INIT_38 => X"42026FC04202586841FFEE4041EC2B7041E6E90041E59E5041E66EB041E3ED30",
--INIT_39 => X"4202E478420578104202DBC842061EF04204D1604209A49842055EF84206CC80",
--INIT_3a => X"41E2030041E6BB3041E5808041E7F58041E73B7041F5551041F6478042021388",
--INIT_3b => X"41E312D041E71A7041E422E041E604C041E437D041E513A041E4998041E46270",
--INIT_3c => X"420361004202B92841F1B20041FCBC0041E810D041E83E3041E3A52041E37060",
--INIT_3d => X"4202FF1042025670420466484203D31842070EA84202FDD04205B4884202FCD8",
--INIT_3e => X"41E2171041E6030041E72CC041E439D041EAD52041E7575042024CB841FAFBE0",
--INIT_3f => X"41E73B3041E5BE4041E4134041E6E52041E3111041E6E8E041E2E42041E38C60",
--INIT_40 => X"420255B84204AFE841FB288041F79C0041EC08E041ED2C8041EDDFB041E99860",
--INIT_41 => X"42016768420653284205AEE8420587904204BB00420711A84204E9D042057EC8",
--INIT_42 => X"41E7F9A041ED55F041E8B91041EA99B041E9178041F1CA6041F15C404204CCC8",
--INIT_43 => X"41F0EE6041EF975041EFCD0041F1866041F21EA041EC0F0041E9D92041E851C0",
--INIT_44 => X"42013C5041F7D7C041F41E1041EC3BA041E88C8041E5DA2041E2A9D041E1BE30",
--INIT_45 => X"4202FAF041FED2C04203AC38420274F842018368420195D04201425841FEED40",
--INIT_46 => X"41E43B6041E1772041E36C9041E5A22041E5A45041E3C97041F91B0041F0FD00",
--INIT_47 => X"41E8174041E6683041EE368041F2B3B041E6232041EBA9F041E5F06041E4C4E0",
--INIT_48 => X"41EB899041EF415041E62F8041E9ED5041E35F6041E52EB041E4A5B041E3FC60",
--INIT_49 => X"41F114E04202A4D8420149D04201581841FF5F904201CB6041F67A2041FDF1F0",
--INIT_4a => X"41E2B1C041E4C07041E563D041E568A041E42CC041EA6D8041E7506041FA0890",
--INIT_4b => X"41EEA83041FCC9504201595041FA12B041FA448041EA676041E62EA041E851C0",
--INIT_4c => X"41EE392041E6929041E511C041E412D041E44AF041E27FA041E1A52041E74D00",
--INIT_4d => X"4200483041F484D042003A3841FDA4B041FD5E1041F3EBA041F443B041EB5F50",
--INIT_4e => X"41E6289041E3064041E267F041E49F3041E46FF041E1FAA041EDA01041E7A270",
--INIT_4f => X"4200D2284201F1F042025AF842034E7841EF234041F7106041E6321041E8B070",
--INIT_50 => X"41E57E8041E3A23041E3552041E5E5F041E3BF0041E2B0C041E4275041E44620",
--INIT_51 => X"41EA367041FA89A041F1C7D041F8980041ECF31041EF027041E663A041EA71B0",
--INIT_52 => X"41E3A24041E43D7041E5024041E4ED4041E4770041E4C1D041E1840041ED4300",
--INIT_53 => X"42001B08420913D0420808984201DCE042015A3841F5523041EE498041E5C6E0",
--INIT_54 => X"41E4BBB041E3D30041E20B3041E51E5041E12DE041E35FF041E310C041E798D0",
--INIT_55 => X"41F2A14041E752D041F3B78041E8AC7041E8A69041E7F40041E55A3041E6FB10",
--INIT_56 => X"41E293D041E2F22041E5173041E5A8E041E2FB9041E217E041E695F041E6AA20",
--INIT_57 => X"4204F3A84202D5D8420522B04207679841FB0C7041FD813041E5441041EF7D00",
--INIT_58 => X"41E2325041E754B041E3EBB041E44C0041E0734041E30DE041E2181041E49400",
--INIT_59 => X"41E3FA9041E8736041E4CA6041E780B041E3B2B041E4549041E359D041E5BFB0",
--INIT_5a => X"41E6D74041E7482041E3337041E2E64041E3206041E7478041E4351041E8F640",
--INIT_5b => X"41F2727042040C184204F0C0420489D84202093041FFEEA041FA2CA041E902E0",
--INIT_5c => X"41E2E84041E339E041E33E3041E38C8041E27DC041E2B24041E1A86041E24AF0",
--INIT_5d => X"41E7ED5041E3531041E575B041E4284041E2D59041E599D041E1573041E26D60",
--INIT_5e => X"41E3C43041E49A4041E3A45041E4539041E1F68041DFFAB041E4A1F041E522F0",
--INIT_5f => X"42001DA841F8CEF04202320842045B1842028E00420280C041F1B11041FD3C00"
--)
GENERIC MAP ( -- XXX image raw
INIT_00 => X"C2E14588C2D2D03CC2D648F4C2D6974CC2BCC362C2BDAD43C2BC6645A5258048",
INIT_01 => X"C30C1700C2F9DFFDC30B93C3C307A67FC30499B0C2F56912C3010AA3C2FA7306",
INIT_02 => X"C2D68548C2CE53ADC2DB1641C2D4872BC2FD120FC2F0F104C2FBE2D8C306CBAB",
INIT_03 => X"C22D5420C229BA68C265ED0BC2843817C29B4151C2954CDFC2B477D8C2AD0D45",
INIT_04 => X"C2F206BBC2E5A83EC2D546A8C2D4CD7AC2C48177C2C03C96C2A66E47C29DEC36",
INIT_05 => X"C3070663C315BDC5C3108669C301CB46C3097E04C3093F65C3062A59C30148CD",
INIT_06 => X"C2C4F5F5C2D7FE2EC2DAE749C3005E50C2F359B0C2FAFDB2C307CF08C30ECEF1",
INIT_07 => X"C237ED08C24BC6CAC280AB08C28B5F56C29CDDB5C2A60C08C2B4C983C2C55354",
INIT_08 => X"C3057B7AC306B1A0C2DF4D37C2EC23B9C2D9D1F3C2CBB904C2B64C82C2B9FAC7",
INIT_09 => X"C30D67F5C31720AFC3136DA3C3127EEAC312363FC309B754C3069E2FC30BAFF6",
INIT_0a => X"C2F0857DC2EC3EFAC3022236C2F1D202C30E0A2AC30F8392C312495BC30C8B16",
INIT_0b => X"C2709ABBC27A5B3DC293B27BC29813AFC2B5078DC2B1EAC4C2D0AED6C2D4A553",
INIT_0c => X"C2F66793C303257FC2F9EC53C2F3484DC2D8D991C2D45E11C2C77B79C2BFAB4B",
INIT_0d => X"C30CEF15C315879FC31D6631C315DAFEC316DB0FC30D0287C30B8742C311AD6E",
INIT_0e => X"C2F0643EC2EC4F63C2F2E7C0C306D282C3079FCDC31472C1C3133945C3155FB0",
INIT_0f => X"C258EA83C28AAF62C29AA4B9C2A661E4C2B4EE40C2C29851C2C7DFFFC2DBD471",
INIT_10 => X"C30A88F6C30887E6C2FC3D4BC3067395C2E1FC28C2D1D37BC2CF97CEC2D115D1",
INIT_11 => X"C326D016C312A675C31D7E0DC31D6C6EC317147AC318F79AC30BADD3C30DB53B",
INIT_12 => X"C3018334C3023770C30418D6C316C78FC30F22BCC318E0D6C31D665BC31D2B1F",
INIT_13 => X"C29C52E4C28402F4C2A295C0C2B236CAC2C8ECD1C2B93514C2F0F87CC2EFDA41",
INIT_14 => X"C3091429C2FE8438C30348C6C304A4F3C2F1CAAFC2E29608C2D74F4AC2D6988E",
INIT_15 => X"C31C9277C32728F3C31C7497C3225C3BC310AE36C30D236AC315EE06C2EEA3AD",
INIT_16 => X"C3009C12C30669F9C3079B3CC35274D9C308A78EC3180DA5C31D6631C3151915",
INIT_17 => X"C28F4B0BC2983D86C2AB1190C2B8F2F6C2C0F91CC2C93AD4C2EE70D9C2F8E53E",
INIT_18 => X"C3049B53C30A6F05C307E343C3047F72C2F312ABC2F688A1C2E0BC32C2DB2616",
INIT_19 => X"C32211A0C3252260C3191130C31C144CC2ECA95EC304F28FC2A1184DC2FD9B2C",
INIT_1a => X"C3093D9CC2FFC986C31BB111C318316BC321CA5BC3188BDBC327EA43C3226475",
INIT_1b => X"C2B10557C2919DAFC2C28585C2C6FE09C2CFB8F7C2E3B992C2F75967C311ECF4",
INIT_1c => X"C311D7FBC309BDA5C3154937C3076431C2FC1CB3C2ED9007C2E021F2C2E095E8",
INIT_1d => X"C31B9469C31E57E9C31C48B7C2FF8E99C2DE4402C29D99E7C2F2ED27C281B78D",
INIT_1e => X"C30E150BC30E90FCC3151A36C3208431C31C52F1C321D27EC3268C60C3259367",
INIT_1f => X"C29FE11BC2ADE071C2B20716C2C1DDEFC2D5D049C2E4C83DC2FE00B3C305EDF4",
INIT_20 => X"C2C4D4CAC30877C0C2FE603DC3108914C2FB9F42C2F132EBC2E23358C2EF92A6",
INIT_21 => X"C309E05AC30C8584C2AAD153C2A36E2CC2635273C2416C19C21EF6E6C2C8BD79",
INIT_22 => X"C30CC603C30EA9ABC32501C4C3191CC5C32297D4C31F9DBEC32645A0C335987C",
INIT_23 => X"C2BDCD73C29CAC12C2C8E0E7C2CA7C55C2E64C02C2E3ACE0C308DDE8C308A2DF",
INIT_24 => X"C3052C34C2BC7D60C30C03D5C302D1E5C309F8B4C3008024C2E8A78CC2E2700A",
INIT_25 => X"C2FA2EB4C2BE45C4C2A5035BC2213AD0C2581AF6C2230B73C2675BDFC2071FBE",
INIT_26 => X"C30B8CFDC3174FE8C3134126C31C52B5C3262C4DC31F9EFCC3237116C317A3FD",
INIT_27 => X"C29CBFBEC2C0734FC2C5F71BC2C6CE0FC2DAB29FC2FD0258C3073905C310A913",
INIT_28 => X"C21D062CC2F7BC01C2EF1CABC3062A28C2F2E638C2F45B96C2DFB5A1C2DDD92A",
INIT_29 => X"C25FCAB3C271B710C225B5D8C22DA021C1F361E3C20618EEC1468E05C241CE81",
INIT_2a => X"C3195ACBC318DD7EC31BECDAC3245162C3229AF0C30A6714C2DF51C3C2E736BF",
INIT_2b => X"C2AB6896C2A5A5D1C2C87AF1C2CCB3FBC2EBCB68C2E4C141C3090CC3C30AC9B5",
INIT_2c => X"C2C20D32C245016BC308D3A1C2E83E3CC2FFC6DAC3066193C2EF3B38C2D8BA9F",
INIT_2d => X"C26FE42EC269A9F4C201BF1CC20D7848C1AB279CC15B1FEDC19B33D541053414",
INIT_2e => X"C30E88DBC3280810C31E9585C327B1B7C311B78DC303720BC2C36F3AC28A4A95",
INIT_2f => X"C29F8C9CC2A5F2EEC2C747ACC2D04ED1C2DDE6F2C2F4234EC30819B0C3177039",
INIT_30 => X"C1411293C2AE48E5C29C7247C3022344C302773FC30ADAD6C2F1E96EC2E68BC6",
INIT_31 => X"C24B3DF4C2329D37C225B5D8C185D649C043EB1740A946B5419455A8C12B767F",
INIT_32 => X"C31461C6C312771AC31D3ABCC3162846C319E464C2AE282DC293FFFAC25D741A",
INIT_33 => X"C2A2C94BC2A7C0ADC2D01BA6C2D3F1BFC2EA4FCCC2F38B04C30F776CC30F489F",
INIT_34 => X"C23195B9C218EC4DC2FD10DDC2AB8B07C3058CFCC2FDDD92C2EB516DC2D6AC95",
INIT_35 => X"C22DA32FC226A2B0C1780B96C190CF5B4184F3C0C021D2E740CBA1C2C02CE22E",
INIT_36 => X"C31C2937C3174A4CC31A65D9C31D4373C2CC0F95C3106CBBC22B9C57C293AB59",
INIT_37 => X"C29E8770C2ABDD87C2BD2B43C2C847FEC2E5A71FC2F8BA3FC308C569C30C1097",
INIT_38 => X"C2156B95C2210246C256AEB5C2EF1CCBC2F1DAE4C2EF71A6C2DC674EC2E352BF",
INIT_39 => X"C21D2151C1AD4E58C21EB340C1832F75C1B5D9A4413138DAC194706CC1255540",
INIT_3a => X"C318082FC30CECBAC319FB79C312AE2FC31883AEC2C9BAFAC2C4ECF2C242B85F",
INIT_3b => X"C2A16683C29CA8CCC2C77D54C2CC0266C2DC6F8BC2E86129C301876AC30766AB",
INIT_3c => X"C1EC3D1CC214D893C2C887FBC28256BCC2E985FFC2E11CA7C2E7F576C2E4372D",
INIT_3d => X"C214767BC237562CC1CF1212C2072768C08B09CCC21E88DEC167BD1AC21663E9",
INIT_3e => X"C3166467C30FF0D7C3126A00C320872CC30A533FC317A9DBC2267482C2A7E7E4",
INIT_3f => X"C28F5B91C2A081F3C2C52AA4C2C65DAFC2DFA669C2DD7DBCC3046931C3087CBB",
INIT_40 => X"C20A4D2BC1B87D56C27DBF16C29671C2C2BFD08FC2B84D87C2A50801C2B32F02",
INIT_41 => X"C23C9EBFC161D35CC17D12FDC1A16E2BC1B365D4C109E7A7C1A58FD8C19B5188",
INIT_42 => X"C2EEF709C2DF0E82C30378C8C303EF61C3054FC0C2D5C727C2DBB3BBC1CE6AC8",
INIT_43 => X"C2460449C25F80F1C283D26DC286A46CC28F5B17C2B1EC95C2D6553EC2E6B1FD",
INIT_44 => X"C227FF58C2A2D886C2AE8454C2DF91C4C2D8A7ADC2E47519C2E184BDC2DC0F60",
INIT_45 => X"C20E6FE4C2844042C1F15170C22F2BCAC237C58EC2448A20C23BA876C27C025B",
INIT_46 => X"C305D929C31796D4C319DE0DC31971D3C3146230C31F56B7C2A73B63C2F15E13",
INIT_47 => X"C283228AC2933AD1C28CEB85C2854F60C2CDDF42C2B94994C2F1CE26C300F237",
INIT_48 => X"C2E4436CC2D84386C2FDB76CC2EF878BC2EEA63BC2E836D7C2D1143DC2CDA36F",
INIT_49 => X"C2DD9EFAC2243C91C247CA49C250BF28C26634D9C235673CC2B590A4C283F5D3",
INIT_4a => X"C305A6ADC305356EC30DCD3AC3141E9EC314814FC305C3E8C314D9E5C2A5D3A8",
INIT_4b => X"C247A2B9C2085697C1D3A210C239B56DC2470DA5C2B8A185C2E4A155C2E6B1FD",
INIT_4c => X"C2D08499C3064C08C2FFCBDEC3073515C2E329CFC2F248C0C2D9AF54C2BC1AB8",
INIT_4d => X"C2572AEFC2C9DA2DC260E13FC28D0191C27D26BAC2C4CE46C2C0E145C3025238",
INIT_4e => X"C2F30AF6C3078FF1C3153059C3147C93C31219D8C321E74DC2F9B066C3147D18",
INIT_4f => X"C19E6A39C1A87939C1A5E0CDC19EBF0DC29189F9C2735B51C2DF1F53C2E0B061",
INIT_50 => X"C2F89F28C3008F7BC2FE8D27C2EE82F8C2DC67A2C2D979A8C2BD5552C2BB625D",
INIT_51 => X"C2FF6EE0C29577DAC2CCE5E9C2A26F6EC2E9C69CC2D6AE36C307E9DEC2F483D2",
INIT_52 => X"C2EA8947C2F7317AC30245DCC308062CC30A850BC310271FC321EFD3C2F4A6B3",
INIT_53 => X"C1AB00604000D18C3F8A2AFAC1CA258AC1D8543FC26F9A37C2A2E8B0C2DC68E2",
INIT_54 => X"C2F6031EC2FAD167C2FE5724C2EC0E51C2E21FFCC2D16B96C2BC9310C2A90B1B",
INIT_55 => X"C2C2CCAEC3091D1EC2BB6C26C303EC77C3002839C300B36AC308C799C303A0CF",
INIT_56 => X"C2EA9F48C2F8E899C2FE3C9FC3025F67C30C334EC31677E4C30CC18AC30F1DE4",
INIT_57 => X"C0CFDA6BC18018AAC100B6A6C03EDBF2C22312A7C2243FB3C2C78742C2A721F9",
INIT_58 => X"C2F5F547C2DD5437C2DBA9FBC2DBBF93C2CCCECCC2C74AEAC2B392ABC2ABFD8C",
INIT_59 => X"C3089B10C2FD8B6AC30AEF89C3062530C2FEE3D4C3056414C30080ABC2FFDF06",
INIT_5a => X"C2C409F4C2CE49E5C2F8871FC3013AF1C2FA1F8CC2F30AE5C308AA36C2FF0A9A",
INIT_5b => X"C20B91DEC13B173AC112EFAFC155D730C1AB0A56C200F7DCC2425A67C2B4C186",
INIT_5c => X"C2E97EC5C2ED9DF5C2D8CE68C2DB9069C2BE8590C2C55A4EC2AF832EC2B1154A",
INIT_5d => X"C2F1835DC30BC15CC304C4AAC30DE924C2FC1A05C2FCD12DC302D9BCC3076A74",
INIT_5e => X"C2CBACB8C2D68459C2ED4372C2F416FFC2F90ED5C30C4E3CC302B874C308C2F0",
INIT_5f => X"C185B163C1F27A56C183F057C15100ABC18CA655C1ADDD82C28219C9C22E807E"
)
PORT MAP (
DO => o_do,
DOP => open,
ADDR => i_addr,
CLK => i_clock,
DI => (others => '0'),
DIP => (others => '0'),
EN => '1',
SSR => i_reset,
WE => '0'
);

end Behavioral;

