----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:57:15 02/07/2023 
-- Design Name: 
-- Module Name:    ExtractOffsetParameters - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE,ieee_proposed;
use IEEE.STD_LOGIC_1164.ALL;

use ieee_proposed.fixed_pkg.all;

USE work.p_fphdl_package1.all;
USE work.p_fphdl_package3.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ExtractOffsetParameters is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_run : in std_logic;

--i_ee0x2410 : in slv16; -- 1-occremscale,2-occcolumnscale,3-occrowscale
--i_offsetRef : in fd2ft; -- offsetref from fixed2float
--
--i_ee0x2412 : in slv16; -- occrow1-4
--i_ee0x2413 : in slv16; -- occrow5-8
--i_ee0x2414 : in slv16; -- occrow9-12
--i_ee0x2415 : in slv16; -- occrow13-16
--i_ee0x2416 : in slv16; -- occrow17-20
--i_ee0x2417 : in slv16; -- occrow21-24
--
--i_ee0x2418 : in slv16; -- occcol1-4
--i_ee0x2419 : in slv16; -- occcol5-8
--i_ee0x241a : in slv16; -- occcol9-12
--i_ee0x241b : in slv16; -- occcol13-16
--i_ee0x241c : in slv16; -- occcol17-20
--i_ee0x241d : in slv16; -- occcol21-24
--i_ee0x241e : in slv16; -- occcol25-28
--i_ee0x241f : in slv16; -- occcol29-32
--
--i_ee0x2440 : in slv16; -- offset ROWS*COLS

i2c_mem_ena : out STD_LOGIC;
i2c_mem_addra : out STD_LOGIC_VECTOR(11 DOWNTO 0);
i2c_mem_douta : in STD_LOGIC_VECTOR(7 DOWNTO 0);

o_do : out std_logic_vector (31 downto 0);
i_addr : in std_logic_vector (9 downto 0); -- 10bit-1024

o_done : out std_logic;
o_rdy : out std_logic
);
end ExtractOffsetParameters;

architecture Behavioral of ExtractOffsetParameters is

COMPONENT fixed2float
PORT (
a : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
operation_nd : IN STD_LOGIC;
clk : IN STD_LOGIC;
sclr : IN STD_LOGIC;
ce : IN STD_LOGIC;
result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
rdy : OUT STD_LOGIC
);
END COMPONENT;

signal fixed2floata : STD_LOGIC_VECTOR(63 DOWNTO 0);
signal fixed2floatond : STD_LOGIC;
signal fixed2floatclk : STD_LOGIC;
signal fixed2floatsclr : STD_LOGIC;
signal fixed2floatce : STD_LOGIC;
signal fixed2floatr : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal fixed2floatrdy : STD_LOGIC;

COMPONENT mulfp
PORT (
a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
operation_nd : IN STD_LOGIC;
clk : IN STD_LOGIC;
sclr : IN STD_LOGIC;
ce : IN STD_LOGIC;
result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
rdy : OUT STD_LOGIC
);
END COMPONENT;

signal mulfpa : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal mulfpb : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal mulfpond : STD_LOGIC;
signal mulfpclk : STD_LOGIC;
signal mulfpsclr : STD_LOGIC;
signal mulfpce : STD_LOGIC;
signal mulfpr : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal mulfprdy : STD_LOGIC;

COMPONENT addfp
PORT (
a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
b : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
operation_nd : IN STD_LOGIC;
clk : IN STD_LOGIC;
sclr : IN STD_LOGIC;
ce : IN STD_LOGIC;
result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
rdy : OUT STD_LOGIC
);
END COMPONENT;

signal addfpa : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal addfpb : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal addfpond : STD_LOGIC;
signal addfpclk : STD_LOGIC;
signal addfpsclr : STD_LOGIC;
signal addfpce : STD_LOGIC;
signal addfpr : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal addfprdy : STD_LOGIC;

component mem_ramb16_s36_x2 is
generic (
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0a : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0b : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0c : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0d : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0e : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0f : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
);
port (
signal DO : out std_logic_vector (31 downto 0);
signal DOP : out std_logic_vector (3 downto 0);
signal ADDR : in std_logic_vector (9 downto 0); -- 10bit-1024
signal CLK : in std_logic;
signal DI : in std_logic_vector (31 downto 0);
signal DIP : in std_logic_vector (3 downto 0);
signal EN : in std_logic;
signal SSR : in std_logic;
signal WE : in std_logic
);
end component mem_ramb16_s36_x2;

signal addra,mux_addr : std_logic_vector (9 downto 0);
signal doa,dia,mux_dia : std_logic_vector (31 downto 0);

signal ena_mux1 : std_logic;

-- xxx nibbles must out in next clock xyxle
signal nibble1,nibble2,nibble4 : std_logic_vector (3 downto 0);
signal nibble3 : std_logic_vector (5 downto 0);
signal out_nibble1,out_nibble2,out_nibble3,out_nibble4 : std_logic_vector (31 downto 0);

signal write_enable : std_logic;

signal rdy : std_logic;

signal stemp1 : std_logic_vector (15 downto 0);

begin

o_rdy <= rdy;
o_do <= doa when rdy = '1' else (others => '0');
mux_addr <= addra when rdy = '0' else i_addr when rdy = '1' else (others => '0');
mux_dia <= dia when rdy = '0' else (others => '0');

p0 : process (i_clock) is
	constant N_COLS : integer := 32;
	constant N_ROWS : integer := 24;
	variable i : integer range 0 to N_ROWS-1;
	variable j : integer range 0 to N_COLS-1;
	variable index : integer range 0 to 15;
	variable k : integer range 0 to N_COLS*N_ROWS-1;
	constant OFFSET_ST : integer := 1665; -- offset start - eeprom max + 1
	constant OFFSET_SZ : integer := N_COLS*N_ROWS; -- offset size
	variable pixgain_index : integer range 0 to OFFSET_SZ - 1;

	type states is (idle,
	occ0,occ1,occ2,occ3,occ4,
	occ5,occ6,occ7,occ8,occ9,
	occ10,occ11,occ12,occ13,occ14,
	occ15,occ16,occ17,occ18,occ19,
	occ20,occ21,occ22,occ23,occ24,
	occ25,occ26,occ27,occ28,occ29,
	occ30,occ31,occ32,occ33,occ34,
	occ35,occ36,occ37,occ38,occ39,
	occ40,occ41,occ42,occ43,occ44,
	occ45,occ46,occ47,occ48,occ49,
	occ50,occ51,occ52,occ53,occ54,
	occ55,occ56,occ57,occ58,occ59,
	
	occ60,occ61,occ62,occ63,occ64,
	occ65,occ66,occ67,occ68,occ69,
	occ70,occ71,occ72,occ73,occ74,
	occ75,occ76,occ77,occ78,occ79,
	occ80,occ81,occ82,occ83,occ84,
	occ85,occ86,occ87,occ88,occ89,
	occ90,occ91,occ92,occ93,occ94,
	occ95,occ96,occ97,occ98,occ99,
	occ100,occ101,occ102,occ103,occ104,
	occ105,occ106,occ107,occ108,occ109,
	
	occ110,occ111,occ112,occ113,occ114,
	occ115,occ116,occ117,occ118,occ119,
	occ120,occ121,occ122,occ123,occ124,
pow0,pow1,pow2,pow3,pow4,pow5,pow6,


s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,

s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,

s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,

s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,

s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,

s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,

s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,

s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,s638,s639,

s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,

s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,s796,s797,s798,s799,

s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,

s880,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,s958,s959,

s960,s961,s962,s963,s964,s965,s966,s967,s968,s969,s970,s971,s972,s973,s974,s975,s976,s977,s978,s979,s980,s981,s982,s983,s984,s985,s986,s987,s988,s989,s990,s991,s992,s993,s994,s995,s996,s997,s998,s999,s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032,s1033,s1034,s1035,s1036,s1037,s1038,s1039,

s1040,s1041,s1042,s1043,s1044,s1045,s1046,s1047,s1048,s1049,s1050,s1051,s1052,s1053,s1054,s1055,s1056,s1057,s1058,s1059,s1060,s1061,s1062,s1063,s1064,s1065,s1066,s1067,s1068,s1069,s1070,s1071,s1072,s1073,s1074,s1075,s1076,s1077,s1078,s1079,s1080,s1081,s1082,s1083,s1084,s1085,s1086,s1087,s1088,s1089,s1090,s1091,s1092,s1093,s1094,s1095,s1096,s1097,s1098,s1099,s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,

s1120,s1121,s1122,s1123,s1124,s1125,s1126,s1127,s1128,s1129,s1130,s1131,s1132,s1133,s1134,s1135,s1136,s1137,s1138,s1139,s1140,s1141,s1142,s1143,s1144,s1145,s1146,s1147,s1148,s1149,s1150,s1151,s1152,s1153,s1154,s1155,s1156,s1157,s1158,s1159,s1160,s1161,s1162,s1163,s1164,s1165,s1166,s1167,s1168,s1169,s1170,s1171,s1172,s1173,s1174,s1175,s1176,s1177,s1178,s1179,s1180,s1181,s1182,s1183,s1184,s1185,s1186,s1187,s1188,s1189,s1190,s1191,s1192,s1193,s1194,s1195,s1196,s1197,s1198,s1199,

s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,s1231,s1232,s1233,s1234,s1235,s1236,s1237,s1238,s1239,s1240,s1241,s1242,s1243,s1244,s1245,s1246,s1247,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255,s1256,s1257,s1258,s1259,s1260,s1261,s1262,s1263,s1264,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272,s1273,s1274,s1275,s1276,s1277,s1278,s1279,

s1280,s1281,s1282,s1283,s1284,s1285,s1286,s1287,s1288,s1289,s1290,s1291,s1292,s1293,s1294,s1295,s1296,s1297,s1298,s1299,s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324,s1325,s1326,s1327,s1328,s1329,s1330,s1331,s1332,s1333,s1334,s1335,s1336,s1337,s1338,s1339,s1340,s1341,s1342,s1343,s1344,s1345,s1346,s1347,s1348,s1349,s1350,s1351,s1352,s1353,s1354,s1355,s1356,s1357,s1358,s1359,

s1360,s1361,s1362,s1363,s1364,s1365,s1366,s1367,s1368,s1369,s1370,s1371,s1372,s1373,s1374,s1375,s1376,s1377,s1378,s1379,s1380,s1381,s1382,s1383,s1384,s1385,s1386,s1387,s1388,s1389,s1390,s1391,s1392,s1393,s1394,s1395,s1396,s1397,s1398,s1399,s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425,s1426,s1427,s1428,s1429,s1430,s1431,s1432,s1433,s1434,s1435,s1436,s1437,s1438,s1439,

s1440,s1441,s1442,s1443,s1444,s1445,s1446,s1447,s1448,s1449,s1450,s1451,s1452,s1453,s1454,s1455,s1456,s1457,s1458,s1459,s1460,s1461,s1462,s1463,s1464,s1465,s1466,s1467,s1468,s1469,s1470,s1471,s1472,s1473,s1474,s1475,s1476,s1477,s1478,s1479,s1480,s1481,s1482,s1483,s1484,s1485,s1486,s1487,s1488,s1489,s1490,s1491,s1492,s1493,s1494,s1495,s1496,s1497,s1498,s1499,s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,

s1520,s1521,s1522,s1523,s1524,s1525,s1526,s1527,s1528,s1529,s1530,s1531,s1532,s1533,s1534,s1535,s1536,s1537,s1538,s1539,s1540,s1541,s1542,s1543,s1544,s1545,s1546,s1547,s1548,s1549,s1550,s1551,s1552,s1553,s1554,s1555,s1556,s1557,s1558,s1559,s1560,s1561,s1562,s1563,s1564,s1565,s1566,s1567,s1568,s1569,s1570,s1571,s1572,s1573,s1574,s1575,s1576,s1577,s1578,s1579,s1580,s1581,s1582,s1583,s1584,s1585,s1586,s1587,s1588,s1589,s1590,s1591,s1592,s1593,s1594,s1595,s1596,s1597,s1598,s1599,

s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624,s1625,s1626,s1627,s1628,s1629,s1630,s1631,s1632,s1633,s1634,s1635,s1636,s1637,s1638,s1639,s1640,s1641,s1642,s1643,s1644,s1645,s1646,s1647,s1648,s1649,s1650,s1651,s1652,s1653,s1654,s1655,s1656,s1657,s1658,s1659,s1660,s1661,s1662,s1663,s1664,s1665,s1666,s1667,s1668,s1669,s1670,s1671,s1672,s1673,s1674,s1675,s1676,s1677,s1678,s1679,

s1680,s1681,s1682,s1683,s1684,s1685,s1686,s1687,s1688,s1689,s1690,s1691,s1692,s1693,s1694,s1695,s1696,s1697,s1698,s1699,s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724,s1725,s1726,s1727,s1728,s1729,s1730,s1731,s1732,s1733,s1734,s1735,s1736,s1737,s1738,s1739,s1740,s1741,s1742,s1743,s1744,s1745,s1746,s1747,s1748,s1749,s1750,s1751,s1752,s1753,s1754,s1755,s1756,s1757,s1758,s1759,

s1760,s1761,s1762,s1763,s1764,s1765,s1766,s1767,s1768,s1769,s1770,s1771,s1772,s1773,s1774,s1775,s1776,s1777,s1778,s1779,s1780,s1781,s1782,s1783,s1784,s1785,s1786,s1787,s1788,s1789,s1790,s1791,s1792,s1793,s1794,s1795,s1796,s1797,s1798,s1799,s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824,s1825,s1826,s1827,s1828,s1829,s1830,s1831,s1832,s1833,s1834,s1835,s1836,s1837,s1838,s1839,

s1840,s1841,s1842,s1843,s1844,s1845,s1846,s1847,s1848,s1849,s1850,s1851,s1852,s1853,s1854,s1855,s1856,s1857,s1858,s1859,s1860,s1861,s1862,s1863,s1864,s1865,s1866,s1867,s1868,s1869,s1870,s1871,s1872,s1873,s1874,s1875,s1876,s1877,s1878,s1879,s1880,s1881,s1882,s1883,s1884,s1885,s1886,s1887,s1888,s1889,s1890,s1891,s1892,s1893,s1894,s1895,s1896,s1897,s1898,s1899,s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,

s1920,s1921,s1922,s1923,s1924,s1925,s1926,s1927,s1928,s1929,s1930,s1931,s1932,s1933,s1934,s1935,s1936,s1937,s1938,s1939,s1940,s1941,s1942,s1943,s1944,s1945,s1946,s1947,s1948,s1949,s1950,s1951,s1952,s1953,s1954,s1955,s1956,s1957,s1958,s1959,s1960,s1961,s1962,s1963,s1964,s1965,s1966,s1967,s1968,s1969,s1970,s1971,s1972,s1973,s1974,s1975,s1976,s1977,s1978,s1979,s1980,s1981,s1982,s1983,s1984,s1985,s1986,s1987,s1988,s1989,s1990,s1991,s1992,s1993,s1994,s1995,s1996,s1997,s1998,s1999,

s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024,s2025,s2026,s2027,s2028,s2029,s2030,s2031,s2032,s2033,s2034,s2035,s2036,s2037,s2038,s2039,s2040,s2041,s2042,s2043,s2044,s2045,s2046,s2047,s2048,s2049,s2050,s2051,s2052,s2053,s2054,s2055,s2056,s2057,s2058,s2059,s2060,s2061,s2062,s2063,s2064,s2065,s2066,s2067,s2068,s2069,s2070,s2071,s2072,s2073,s2074,s2075,s2076,s2077,s2078,s2079,

s2080,s2081,s2082,s2083,s2084,s2085,s2086,s2087,s2088,s2089,s2090,s2091,s2092,s2093,s2094,s2095,s2096,s2097,s2098,s2099,s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124,s2125,s2126,s2127,s2128,s2129,s2130,s2131,s2132,s2133,s2134,s2135,s2136,s2137,s2138,s2139,s2140,s2141,s2142,s2143,s2144,s2145,s2146,s2147,s2148,s2149,s2150,s2151,s2152,s2153,s2154,s2155,s2156,s2157,s2158,s2159,

s2160,s2161,s2162,s2163,s2164,s2165,s2166,s2167,s2168,s2169,s2170,s2171,s2172,s2173,s2174,s2175,s2176,s2177,s2178,s2179,s2180,s2181,s2182,s2183,s2184,s2185,s2186,s2187,s2188,s2189,s2190,s2191,s2192,s2193,s2194,s2195,s2196,s2197,s2198,s2199,s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224,s2225,s2226,s2227,s2228,s2229,s2230,s2231,s2232,s2233,s2234,s2235,s2236,s2237,s2238,s2239,

s2240,s2241,s2242,s2243,s2244,s2245,s2246,s2247,s2248,s2249,s2250,s2251,s2252,s2253,s2254,s2255,s2256,s2257,s2258,s2259,s2260,s2261,s2262,s2263,s2264,s2265,s2266,s2267,s2268,s2269,s2270,s2271,s2272,s2273,s2274,s2275,s2276,s2277,s2278,s2279,s2280,s2281,s2282,s2283,s2284,s2285,s2286,s2287,s2288,s2289,s2290,s2291,s2292,s2293,s2294,s2295,s2296,s2297,s2298,s2299,s2300,s2301,s2302,s2303,s2304,s2305,s2306,s2307,s2308,s2309,s2310,s2311,s2312,s2313,s2314,s2315,s2316,s2317,s2318,s2319,

s2320,s2321,s2322,s2323,s2324,s2325,s2326,s2327,s2328,s2329,s2330,s2331,s2332,s2333,s2334,s2335,s2336,s2337,s2338,s2339,s2340,s2341,s2342,s2343,s2344,s2345,s2346,s2347,s2348,s2349,s2350,s2351,s2352,s2353,s2354,s2355,s2356,s2357,s2358,s2359,s2360,s2361,s2362,s2363,s2364,s2365,s2366,s2367,s2368,s2369,s2370,s2371,s2372,s2373,s2374,s2375,s2376,s2377,s2378,s2379,s2380,s2381,s2382,s2383,s2384,s2385,s2386,s2387,s2388,s2389,s2390,s2391,s2392,s2393,s2394,s2395,s2396,s2397,s2398,s2399,

s2400,s2401,s2402,s2403,s2404,s2405,s2406,s2407,s2408,s2409,s2410,s2411,s2412,s2413,s2414,s2415,s2416,s2417,s2418,s2419,s2420,s2421,s2422,s2423,s2424,s2425,s2426,s2427,s2428,s2429,s2430,s2431,s2432,s2433,s2434,s2435,s2436,s2437,s2438,s2439,s2440,s2441,s2442,s2443,s2444,s2445,s2446,s2447,s2448,s2449,s2450,s2451,s2452,s2453,s2454,s2455,s2456,s2457,s2458,s2459,s2460,s2461,s2462,s2463,s2464,s2465,s2466,s2467,s2468,s2469,s2470,s2471,s2472,s2473,s2474,s2475,s2476,s2477,s2478,s2479,

s2480,s2481,s2482,s2483,s2484,s2485,s2486,s2487,s2488,s2489,s2490,s2491,s2492,s2493,s2494,s2495,s2496,s2497,s2498,s2499,s2500,s2501,s2502,s2503,s2504,s2505,s2506,s2507,s2508,s2509,s2510,s2511,s2512,s2513,s2514,s2515,s2516,s2517,s2518,s2519,s2520,s2521,s2522,s2523,s2524,s2525,s2526,s2527,s2528,s2529,s2530,s2531,s2532,s2533,s2534,s2535,s2536,s2537,s2538,s2539,s2540,s2541,s2542,s2543,s2544,s2545,s2546,s2547,s2548,s2549,s2550,s2551,s2552,s2553,s2554,s2555,s2556,s2557,s2558,s2559,

s2560,s2561,s2562,s2563,s2564,s2565,s2566,s2567,s2568,s2569,s2570,s2571,s2572,s2573,s2574,s2575,s2576,s2577,s2578,s2579,s2580,s2581,s2582,s2583,s2584,s2585,s2586,s2587,s2588,s2589,s2590,s2591,s2592,s2593,s2594,s2595,s2596,s2597,s2598,s2599,s2600,s2601,s2602,s2603,s2604,s2605,s2606,s2607,s2608,s2609,s2610,s2611,s2612,s2613,s2614,s2615,s2616,s2617,s2618,s2619,s2620,s2621,s2622,s2623,s2624,s2625,s2626,s2627,s2628,s2629,s2630,s2631,s2632,s2633,s2634,s2635,s2636,s2637,s2638,s2639,

s2640,s2641,s2642,s2643,s2644,s2645,s2646,s2647,s2648,s2649,s2650,s2651,s2652,s2653,s2654,s2655,s2656,s2657,s2658,s2659,s2660,s2661,s2662,s2663,s2664,s2665,s2666,s2667,s2668,s2669,s2670,s2671,s2672,s2673,s2674,s2675,s2676,s2677,s2678,s2679,s2680,s2681,s2682,s2683,s2684,s2685,s2686,s2687,s2688,s2689,s2690,s2691,s2692,s2693,s2694,s2695,s2696,s2697,s2698,s2699,s2700,s2701,s2702,s2703,s2704,s2705,s2706,s2707,s2708,s2709,s2710,s2711,s2712,s2713,s2714,s2715,s2716,s2717,s2718,s2719,

s2720,s2721,s2722,s2723,s2724,s2725,s2726,s2727,s2728,s2729,s2730,s2731,s2732,s2733,s2734,s2735,s2736,s2737,s2738,s2739,s2740,s2741,s2742,s2743,s2744,s2745,s2746,s2747,s2748,s2749,s2750,s2751,s2752,s2753,s2754,s2755,s2756,s2757,s2758,s2759,s2760,s2761,s2762,s2763,s2764,s2765,s2766,s2767,s2768,s2769,s2770,s2771,s2772,s2773,s2774,s2775,s2776,s2777,s2778,s2779,s2780,s2781,s2782,s2783,s2784,s2785,s2786,s2787,s2788,s2789,s2790,s2791,s2792,s2793,s2794,s2795,s2796,s2797,s2798,s2799,

s2800,s2801,s2802,s2803,s2804,s2805,s2806,s2807,s2808,s2809,s2810,s2811,s2812,s2813,s2814,s2815,s2816,s2817,s2818,s2819,s2820,s2821,s2822,s2823,s2824,s2825,s2826,s2827,s2828,s2829,s2830,s2831,s2832,s2833,s2834,s2835,s2836,s2837,s2838,s2839,s2840,s2841,s2842,s2843,s2844,s2845,s2846,s2847,s2848,s2849,s2850,s2851,s2852,s2853,s2854,s2855,s2856,s2857,s2858,s2859,s2860,s2861,s2862,s2863,s2864,s2865,s2866,s2867,s2868,s2869,s2870,s2871,s2872,s2873,s2874,s2875,s2876,s2877,s2878,s2879,

s2880,s2881,s2882,s2883,s2884,s2885,s2886,s2887,s2888,s2889,s2890,s2891,s2892,s2893,s2894,s2895,s2896,s2897,s2898,s2899,s2900,s2901,s2902,s2903,s2904,s2905,s2906,s2907,s2908,s2909,s2910,s2911,s2912,s2913,s2914,s2915,s2916,s2917,s2918,s2919,s2920,s2921,s2922,s2923,s2924,s2925,s2926,s2927,s2928,s2929,s2930,s2931,s2932,s2933,s2934,s2935,s2936,s2937,s2938,s2939,s2940,s2941,s2942,s2943,s2944,s2945,s2946,s2947,s2948,s2949,s2950,s2951,s2952,s2953,s2954,s2955,s2956,s2957,s2958,s2959,

s2960,s2961,s2962,s2963,s2964,s2965,s2966,s2967,s2968,s2969,s2970,s2971,s2972,s2973,s2974,s2975,s2976,s2977,s2978,s2979,s2980,s2981,s2982,s2983,s2984,s2985,s2986,s2987,s2988,s2989,s2990,s2991,s2992,s2993,s2994,s2995,s2996,s2997,s2998,s2999,s3000,s3001,s3002,s3003,s3004,s3005,s3006,s3007,s3008,s3009,s3010,s3011,s3012,s3013,s3014,s3015,s3016,s3017,s3018,s3019,s3020,s3021,s3022,s3023,s3024,s3025,s3026,s3027,s3028,s3029,s3030,s3031,s3032,s3033,s3034,s3035,s3036,s3037,s3038,s3039,

s3040,s3041,s3042,s3043,s3044,s3045,s3046,s3047,s3048,s3049,s3050,s3051,s3052,s3053,s3054,s3055,s3056,s3057,s3058,s3059,s3060,s3061,s3062,s3063,s3064,s3065,s3066,s3067,s3068,s3069,s3070,s3071,s3072,s3073,s3074,s3075,s3076,s3077,s3078,s3079,s3080,s3081,s3082,s3083,s3084,s3085,s3086,s3087,s3088,s3089,s3090,s3091,s3092,s3093,s3094,s3095,s3096,s3097,s3098,s3099,s3100,s3101,s3102,s3103,s3104,s3105,s3106,s3107,s3108,s3109,s3110,s3111,s3112,s3113,s3114,s3115,s3116,s3117,s3118,s3119,

s3120,s3121,s3122,s3123,s3124,s3125,s3126,s3127,s3128,s3129,s3130,s3131,s3132,s3133,s3134,s3135,s3136,s3137,s3138,s3139,s3140,s3141,s3142,s3143,s3144,s3145,s3146,s3147,s3148,s3149,s3150,s3151,s3152,s3153,s3154,s3155,s3156,s3157,s3158,s3159,s3160,s3161,s3162,s3163,s3164,s3165,s3166,s3167,s3168,s3169,s3170,s3171,s3172,s3173,s3174,s3175,s3176,s3177,s3178,s3179,s3180,s3181,s3182,s3183,s3184,s3185,s3186,s3187,s3188,s3189,s3190,s3191,s3192,s3193,s3194,s3195,s3196,s3197,s3198,s3199,

s3200,s3201,s3202,s3203,s3204,s3205,s3206,s3207,s3208,s3209,s3210,s3211,s3212,s3213,s3214,s3215,s3216,s3217,s3218,s3219,s3220,s3221,s3222,s3223,s3224,s3225,s3226,s3227,s3228,s3229,s3230,s3231,s3232,s3233,s3234,s3235,s3236,s3237,s3238,s3239,s3240,s3241,s3242,s3243,s3244,s3245,s3246,s3247,s3248,s3249,s3250,s3251,s3252,s3253,s3254,s3255,s3256,s3257,s3258,s3259,s3260,s3261,s3262,s3263,s3264,s3265,s3266,s3267,s3268,s3269,s3270,s3271,s3272,s3273,s3274,s3275,s3276,s3277,s3278,s3279,

s3280,s3281,s3282,s3283,s3284,s3285,s3286,s3287,s3288,s3289,s3290,s3291,s3292,s3293,s3294,s3295,s3296,s3297,s3298,s3299,s3300,s3301,s3302,s3303,s3304,s3305,s3306,s3307,s3308,s3309,s3310,s3311,s3312,s3313,s3314,s3315,s3316,s3317,s3318,s3319,s3320,s3321,s3322,s3323,s3324,s3325,s3326,s3327,s3328,s3329,s3330,s3331,s3332,s3333,s3334,s3335,s3336,s3337,s3338,s3339,s3340,s3341,s3342,s3343,s3344,s3345,s3346,s3347,s3348,s3349,s3350,s3351,s3352,s3353,s3354,s3355,s3356,s3357,s3358,s3359,

s3360,s3361,s3362,s3363,s3364,s3365,s3366,s3367,s3368,s3369,s3370,s3371,s3372,s3373,s3374,s3375,s3376,s3377,s3378,s3379,s3380,s3381,s3382,s3383,s3384,s3385,s3386,s3387,s3388,s3389,s3390,s3391,s3392,s3393,s3394,s3395,s3396,s3397,s3398,s3399,s3400,s3401,s3402,s3403,s3404,s3405,s3406,s3407,s3408,s3409,s3410,s3411,s3412,s3413,s3414,s3415,s3416,s3417,s3418,s3419,s3420,s3421,s3422,s3423,s3424,s3425,s3426,s3427,s3428,s3429,s3430,s3431,s3432,s3433,s3434,s3435,s3436,s3437,s3438,s3439,

s3440,s3441,s3442,s3443,s3444,s3445,s3446,s3447,s3448,s3449,s3450,s3451,s3452,s3453,s3454,s3455,s3456,s3457,s3458,s3459,s3460,s3461,s3462,s3463,s3464,s3465,s3466,s3467,s3468,s3469,s3470,s3471,s3472,s3473,s3474,s3475,s3476,s3477,s3478,s3479,s3480,s3481,s3482,s3483,s3484,s3485,s3486,s3487,s3488,s3489,s3490,s3491,s3492,s3493,s3494,s3495,s3496,s3497,s3498,s3499,s3500,s3501,s3502,s3503,s3504,s3505,s3506,s3507,s3508,s3509,s3510,s3511,s3512,s3513,s3514,s3515,s3516,s3517,s3518,s3519,

s3520,s3521,s3522,s3523,s3524,s3525,s3526,s3527,s3528,s3529,s3530,s3531,s3532,s3533,s3534,s3535,s3536,s3537,s3538,s3539,s3540,s3541,s3542,s3543,s3544,s3545,s3546,s3547,s3548,s3549,s3550,s3551,s3552,s3553,s3554,s3555,s3556,s3557,s3558,s3559,s3560,s3561,s3562,s3563,s3564,s3565,s3566,s3567,s3568,s3569,s3570,s3571,s3572,s3573,s3574,s3575,s3576,s3577,s3578,s3579,s3580,s3581,s3582,s3583,s3584,s3585,s3586,s3587,s3588,s3589,s3590,s3591,s3592,s3593,s3594,s3595,s3596,s3597,s3598,s3599,

s3600,s3601,s3602,s3603,s3604,s3605,s3606,s3607,s3608,s3609,s3610,s3611,s3612,s3613,s3614,s3615,s3616,s3617,s3618,s3619,s3620,s3621,s3622,s3623,s3624,s3625,s3626,s3627,s3628,s3629,s3630,s3631,s3632,s3633,s3634,s3635,s3636,s3637,s3638,s3639,s3640,s3641,s3642,s3643,s3644,s3645,s3646,s3647,s3648,s3649,s3650,s3651,s3652,s3653,s3654,s3655,s3656,s3657,s3658,s3659,s3660,s3661,s3662,s3663,s3664,s3665,s3666,s3667,s3668,s3669,s3670,s3671,s3672,s3673,s3674,s3675,s3676,s3677,s3678,s3679,

s3680,s3681,s3682,s3683,s3684,s3685,s3686,s3687,s3688,s3689,s3690,s3691,s3692,s3693,s3694,s3695,s3696,s3697,s3698,s3699,s3700,s3701,s3702,s3703,s3704,s3705,s3706,s3707,s3708,s3709,s3710,s3711,s3712,s3713,s3714,s3715,s3716,s3717,s3718,s3719,s3720,s3721,s3722,s3723,s3724,s3725,s3726,s3727,s3728,s3729,s3730,s3731,s3732,s3733,s3734,s3735,s3736,s3737,s3738,s3739,s3740,s3741,s3742,s3743,s3744,s3745,s3746,s3747,s3748,s3749,s3750,s3751,s3752,s3753,s3754,s3755,s3756,s3757,s3758,s3759,

s3760,s3761,s3762,s3763,s3764,s3765,s3766,s3767,s3768,s3769,s3770,s3771,s3772,s3773,s3774,s3775,s3776,s3777,s3778,s3779,s3780,s3781,s3782,s3783,s3784,s3785,s3786,s3787,s3788,s3789,s3790,s3791,s3792,s3793,s3794,s3795,s3796,s3797,s3798,s3799,s3800,s3801,s3802,s3803,s3804,s3805,s3806,s3807,s3808,s3809,s3810,s3811,s3812,s3813,s3814,s3815,s3816,s3817,s3818,s3819,s3820,s3821,s3822,s3823,s3824,s3825,s3826,s3827,s3828,s3829,s3830,s3831,s3832,s3833,s3834,s3835,s3836,s3837,s3838,s3839,

s3840,s3841,s3842,s3843,s3844,s3845,s3846,s3847,s3848,s3849,s3850,s3851,s3852,s3853,s3854,s3855,s3856,s3857,s3858,s3859,s3860,s3861,s3862,s3863,s3864,s3865,s3866,s3867,s3868,s3869,s3870,s3871,s3872,s3873,s3874,s3875,s3876,s3877,s3878,s3879,s3880,s3881,s3882,s3883,s3884,s3885,s3886,s3887,s3888,s3889,s3890,s3891,s3892,s3893,s3894,s3895,s3896,s3897,s3898,s3899,s3900,s3901,s3902,s3903,s3904,s3905,s3906,s3907,s3908,s3909,s3910,s3911,s3912,s3913,s3914,s3915,s3916,s3917,s3918,s3919,

s3920,s3921,s3922,s3923,s3924,s3925,s3926,s3927,s3928,s3929,s3930,s3931,s3932,s3933,s3934,s3935,s3936,s3937,s3938,s3939,s3940,s3941,s3942,s3943,s3944,s3945,s3946,s3947,s3948,s3949,s3950,s3951,s3952,s3953,s3954,s3955,s3956,s3957,s3958,s3959,s3960,s3961,s3962,s3963,s3964,s3965,s3966,s3967,s3968,s3969,s3970,s3971,s3972,s3973,s3974,s3975,s3976,s3977,s3978,s3979,s3980,s3981,s3982,s3983,s3984,s3985,s3986,s3987,s3988,s3989,s3990,s3991,s3992,s3993,s3994,s3995,s3996,s3997,s3998,s3999,

s4000,s4001,s4002,s4003,s4004,s4005,s4006,s4007,s4008,s4009,s4010,s4011,s4012,s4013,s4014,s4015,s4016,s4017,s4018,s4019,s4020,s4021,s4022,s4023,s4024,s4025,s4026,s4027,s4028,s4029,s4030,s4031,s4032,s4033,s4034,s4035,s4036,s4037,s4038,s4039,s4040,s4041,s4042,s4043,s4044,s4045,s4046,s4047,s4048,s4049,s4050,s4051,s4052,s4053,s4054,s4055,s4056,s4057,s4058,s4059,s4060,s4061,s4062,s4063,s4064,s4065,s4066,s4067,s4068,s4069,s4070,s4071,s4072,s4073,s4074,s4075,s4076,s4077,s4078,s4079,

s4080,s4081,s4082,s4083,s4084,s4085,s4086,s4087,s4088,s4089,s4090,s4091,s4092,s4093,s4094,s4095,s4096,s4097,s4098,s4099,s4100,s4101,s4102,s4103,s4104,s4105,s4106,s4107,s4108,s4109,s4110,s4111,s4112,s4113,s4114,s4115,s4116,s4117,s4118,s4119,s4120,s4121,s4122,s4123,s4124,s4125,s4126,s4127,s4128,s4129,s4130,s4131,s4132,s4133,s4134,s4135,s4136,s4137,s4138,s4139,s4140,s4141,s4142,s4143,s4144,s4145,s4146,s4147,s4148,s4149,s4150,s4151,s4152,s4153,s4154,s4155,s4156,s4157,s4158,s4159,

s4160,s4161,s4162,s4163,s4164,s4165,s4166,s4167,s4168,s4169,s4170,s4171,s4172,s4173,s4174,s4175,s4176,s4177,s4178,s4179,s4180,s4181,s4182,s4183,s4184,s4185,s4186,s4187,s4188,s4189,s4190,s4191,s4192,s4193,s4194,s4195,s4196,s4197,s4198,s4199,s4200,s4201,s4202,s4203,s4204,s4205,s4206,s4207,s4208,s4209,s4210,s4211,s4212,s4213,s4214,s4215,s4216,s4217,s4218,s4219,s4220,s4221,s4222,s4223,s4224,s4225,s4226,s4227,s4228,s4229,s4230,s4231,s4232,s4233,s4234,s4235,s4236,s4237,s4238,s4239,

s4240,s4241,s4242,s4243,s4244,s4245,s4246,s4247,s4248,s4249,s4250,s4251,s4252,s4253,s4254,s4255,s4256,s4257,s4258,s4259,s4260,s4261,s4262,s4263,s4264,s4265,s4266,s4267,s4268,s4269,s4270,s4271,s4272,s4273,s4274,s4275,s4276,s4277,s4278,s4279,s4280,s4281,s4282,s4283,s4284,s4285,s4286,s4287,s4288,s4289,s4290,s4291,s4292,s4293,s4294,s4295,s4296,s4297,s4298,s4299,s4300,s4301,s4302,s4303,s4304,s4305,s4306,s4307,s4308,s4309,s4310,s4311,s4312,s4313,s4314,s4315,s4316,s4317,s4318,s4319,

s4320,s4321,s4322,s4323,s4324,s4325,s4326,s4327,s4328,s4329,s4330,s4331,s4332,s4333,s4334,s4335,s4336,s4337,s4338,s4339,s4340,s4341,s4342,s4343,s4344,s4345,s4346,s4347,s4348,s4349,s4350,s4351,s4352,s4353,s4354,s4355,s4356,s4357,s4358,s4359,s4360,s4361,s4362,s4363,s4364,s4365,s4366,s4367,s4368,s4369,s4370,s4371,s4372,s4373,s4374,s4375,s4376,s4377,s4378,s4379,s4380,s4381,s4382,s4383,s4384,s4385,s4386,s4387,s4388,s4389,s4390,s4391,s4392,s4393,s4394,s4395,s4396,s4397,s4398,s4399,

s4400,s4401,s4402,s4403,s4404,s4405,s4406,s4407,s4408,s4409,s4410,s4411,s4412,s4413,s4414,s4415,s4416,s4417,s4418,s4419,s4420,s4421,s4422,s4423,s4424,s4425,s4426,s4427,s4428,s4429,s4430,s4431,s4432,s4433,s4434,s4435,s4436,s4437,s4438,s4439,s4440,s4441,s4442,s4443,s4444,s4445,s4446,s4447,s4448,s4449,s4450,s4451,s4452,s4453,s4454,s4455,s4456,s4457,s4458,s4459,s4460,s4461,s4462,s4463,s4464,s4465,s4466,s4467,s4468,s4469,s4470,s4471,s4472,s4473,s4474,s4475,s4476,s4477,s4478,s4479,

s4480,s4481,s4482,s4483,s4484,s4485,s4486,s4487,s4488,s4489,s4490,s4491,s4492,s4493,s4494,s4495,s4496,s4497,s4498,s4499,s4500,s4501,s4502,s4503,s4504,s4505,s4506,s4507,s4508,s4509,s4510,s4511,s4512,s4513,s4514,s4515,s4516,s4517,s4518,s4519,s4520,s4521,s4522,s4523,s4524,s4525,s4526,s4527,s4528,s4529,s4530,s4531,s4532,s4533,s4534,s4535,s4536,s4537,s4538,s4539,s4540,s4541,s4542,s4543,s4544,s4545,s4546,s4547,s4548,s4549,s4550,s4551,s4552,s4553,s4554,s4555,s4556,s4557,s4558,s4559,

s4560,s4561,s4562,s4563,s4564,s4565,s4566,s4567,s4568,s4569,s4570,s4571,s4572,s4573,s4574,s4575,s4576,s4577,s4578,s4579,s4580,s4581,s4582,s4583,s4584,s4585,s4586,s4587,s4588,s4589,s4590,s4591,s4592,s4593,s4594,s4595,s4596,s4597,s4598,s4599,s4600,s4601,s4602,s4603,s4604,s4605,s4606,s4607,s4608,s4609,s4610,s4611,s4612,s4613,s4614,s4615,s4616,s4617,s4618,s4619,s4620,s4621,s4622,s4623,s4624,s4625,s4626,s4627,s4628,s4629,s4630,s4631,s4632,s4633,s4634,s4635,s4636,s4637,s4638,s4639,

s4640,s4641,s4642,s4643,s4644,s4645,s4646,s4647,s4648,s4649,s4650,s4651,s4652,s4653,s4654,s4655,s4656,s4657,s4658,s4659,s4660,s4661,s4662,s4663,s4664,s4665,s4666,s4667,s4668,s4669,s4670,s4671,s4672,s4673,s4674,s4675,s4676,s4677,s4678,s4679,s4680,s4681,s4682,s4683,s4684,s4685,s4686,s4687,s4688,s4689,s4690,s4691,s4692,s4693,s4694,s4695,s4696,s4697,s4698,s4699,s4700,s4701,s4702,s4703,s4704,s4705,s4706,s4707,s4708,s4709,s4710,s4711,s4712,s4713,s4714,s4715,s4716,s4717,s4718,s4719,

s4720,s4721,s4722,s4723,s4724,s4725,s4726,s4727,s4728,s4729,s4730,s4731,s4732,s4733,s4734,s4735,s4736,s4737,s4738,s4739,s4740,s4741,s4742,s4743,s4744,s4745,s4746,s4747,s4748,s4749,s4750,s4751,s4752,s4753,s4754,s4755,s4756,s4757,s4758,s4759,s4760,s4761,s4762,s4763,s4764,s4765,s4766,s4767,s4768,s4769,s4770,s4771,s4772,s4773,s4774,s4775,s4776,s4777,s4778,s4779,s4780,s4781,s4782,s4783,s4784,s4785,s4786,s4787,s4788,s4789,s4790,s4791,s4792,s4793,s4794,s4795,s4796,s4797,s4798,s4799,

s4800,s4801,s4802,s4803,s4804,s4805,s4806,s4807,s4808,s4809,s4810,s4811,s4812,s4813,s4814,s4815,s4816,s4817,s4818,s4819,s4820,s4821,s4822,s4823,s4824,s4825,s4826,s4827,s4828,s4829,s4830,s4831,s4832,s4833,s4834,s4835,s4836,s4837,s4838,s4839,s4840,s4841,s4842,s4843,s4844,s4845,s4846,s4847,s4848,s4849,s4850,s4851,s4852,s4853,s4854,s4855,s4856,s4857,s4858,s4859,s4860,s4861,s4862,s4863,s4864,s4865,s4866,s4867,s4868,s4869,s4870,s4871,s4872,s4873,s4874,s4875,s4876,s4877,s4878,s4879,

s4880,s4881,s4882,s4883,s4884,s4885,s4886,s4887,s4888,s4889,s4890,s4891,s4892,s4893,s4894,s4895,s4896,s4897,s4898,s4899,s4900,s4901,s4902,s4903,s4904,s4905,s4906,s4907,s4908,s4909,s4910,s4911,s4912,s4913,s4914,s4915,s4916,s4917,s4918,s4919,s4920,s4921,s4922,s4923,s4924,s4925,s4926,s4927,s4928,s4929,s4930,s4931,s4932,s4933,s4934,s4935,s4936,s4937,s4938,s4939,s4940,s4941,s4942,s4943,s4944,s4945,s4946,s4947,s4948,s4949,s4950,s4951,s4952,s4953,s4954,s4955,s4956,s4957,s4958,s4959,

s4960,s4961,s4962,s4963,s4964,s4965,s4966,s4967,s4968,s4969,s4970,s4971,s4972,s4973,s4974,s4975,s4976,s4977,s4978,s4979,s4980,s4981,s4982,s4983,s4984,s4985,s4986,s4987,s4988,s4989,s4990,s4991,s4992,s4993,s4994,s4995,s4996,s4997,s4998,s4999,s5000,s5001,s5002,s5003,s5004,s5005,s5006,s5007,s5008,s5009,s5010,s5011,s5012,s5013,s5014,s5015,s5016,s5017,s5018,s5019,s5020,s5021,s5022,s5023,s5024,s5025,s5026,s5027,s5028,s5029,s5030,s5031,s5032,s5033,s5034,s5035,s5036,s5037,s5038,s5039,

s5040,s5041,s5042,s5043,s5044,s5045,s5046,s5047,s5048,s5049,s5050,s5051,s5052,s5053,s5054,s5055,s5056,s5057,s5058,s5059,s5060,s5061,s5062,s5063,s5064,s5065,s5066,s5067,s5068,s5069,s5070,s5071,s5072,s5073,s5074,s5075,s5076,s5077,s5078,s5079,s5080,s5081,s5082,s5083,s5084,s5085,s5086,s5087,s5088,s5089,s5090,s5091,s5092,s5093,s5094,s5095,s5096,s5097,s5098,s5099,s5100,s5101,s5102,s5103,s5104,s5105,s5106,s5107,s5108,s5109,s5110,s5111,s5112,s5113,s5114,s5115,s5116,s5117,s5118,s5119,

s5120,s5121,s5122,s5123,s5124,s5125,s5126,s5127,s5128,s5129,s5130,s5131,s5132,s5133,s5134,s5135,s5136,s5137,s5138,s5139,s5140,s5141,s5142,s5143,s5144,s5145,s5146,s5147,s5148,s5149,s5150,s5151,s5152,s5153,s5154,s5155,s5156,s5157,s5158,s5159,s5160,s5161,s5162,s5163,s5164,s5165,s5166,s5167,s5168,s5169,s5170,s5171,s5172,s5173,s5174,s5175,s5176,s5177,s5178,s5179,s5180,s5181,s5182,s5183,s5184,s5185,s5186,s5187,s5188,s5189,s5190,s5191,s5192,s5193,s5194,s5195,s5196,s5197,s5198,s5199,

s5200,s5201,s5202,s5203,s5204,s5205,s5206,s5207,s5208,s5209,s5210,s5211,s5212,s5213,s5214,s5215,s5216,s5217,s5218,s5219,s5220,s5221,s5222,s5223,s5224,s5225,s5226,s5227,s5228,s5229,s5230,s5231,s5232,s5233,s5234,s5235,s5236,s5237,s5238,s5239,s5240,s5241,s5242,s5243,s5244,s5245,s5246,s5247,s5248,s5249,s5250,s5251,s5252,s5253,s5254,s5255,s5256,s5257,s5258,s5259,s5260,s5261,s5262,s5263,s5264,s5265,s5266,s5267,s5268,s5269,s5270,s5271,s5272,s5273,s5274,s5275,s5276,s5277,s5278,s5279,

s5280,s5281,s5282,s5283,s5284,s5285,s5286,s5287,s5288,s5289,s5290,s5291,s5292,s5293,s5294,s5295,s5296,s5297,s5298,s5299,s5300,s5301,s5302,s5303,s5304,s5305,s5306,s5307,s5308,s5309,s5310,s5311,s5312,s5313,s5314,s5315,s5316,s5317,s5318,s5319,s5320,s5321,s5322,s5323,s5324,s5325,s5326,s5327,s5328,s5329,s5330,s5331,s5332,s5333,s5334,s5335,s5336,s5337,s5338,s5339,s5340,s5341,s5342,s5343,s5344,s5345,s5346,s5347,s5348,s5349,s5350,s5351,s5352,s5353,s5354,s5355,s5356,s5357,s5358,s5359,

s5360,s5361,s5362,s5363,s5364,s5365,s5366,s5367,s5368,s5369,s5370,s5371,s5372,s5373,s5374,s5375,s5376,s5377,s5378,s5379,s5380,s5381,s5382,s5383,s5384,s5385,s5386,s5387,s5388,s5389,s5390,s5391,s5392,s5393,s5394,s5395,s5396,s5397,s5398,s5399,s5400,s5401,s5402,s5403,s5404,s5405,s5406,s5407,s5408,s5409,s5410,s5411,s5412,s5413,s5414,s5415,s5416,s5417,s5418,s5419,s5420,s5421,s5422,s5423,s5424,s5425,s5426,s5427,s5428,s5429,s5430,s5431,s5432,s5433,s5434,s5435,s5436,s5437,s5438,s5439,

s5440,s5441,s5442,s5443,s5444,s5445,s5446,s5447,s5448,s5449,s5450,s5451,s5452,s5453,s5454,s5455,s5456,s5457,s5458,s5459,s5460,s5461,s5462,s5463,s5464,s5465,s5466,s5467,s5468,s5469,s5470,s5471,s5472,s5473,s5474,s5475,s5476,s5477,s5478,s5479,s5480,s5481,s5482,s5483,s5484,s5485,s5486,s5487,s5488,s5489,s5490,s5491,s5492,s5493,s5494,s5495,s5496,s5497,s5498,s5499,s5500,s5501,s5502,s5503,s5504,s5505,s5506,s5507,s5508,s5509,s5510,s5511,s5512,s5513,s5514,s5515,s5516,s5517,s5518,s5519,

s5520,s5521,s5522,s5523,s5524,s5525,s5526,s5527,s5528,s5529,s5530,s5531,s5532,s5533,s5534,s5535,s5536,s5537,s5538,s5539,s5540,s5541,s5542,s5543,s5544,s5545,s5546,s5547,s5548,s5549,s5550,s5551,s5552,s5553,s5554,s5555,s5556,s5557,s5558,s5559,s5560,s5561,s5562,s5563,s5564,s5565,s5566,s5567,s5568,s5569,s5570,s5571,s5572,s5573,s5574,s5575,s5576,s5577,s5578,s5579,s5580,s5581,s5582,s5583,s5584,s5585,s5586,s5587,s5588,s5589,s5590,s5591,s5592,s5593,s5594,s5595,s5596,s5597,s5598,s5599,

s5600,s5601,s5602,s5603,s5604,s5605,s5606,s5607,s5608,s5609,s5610,s5611,s5612,s5613,s5614,s5615,s5616,s5617,s5618,s5619,s5620,s5621,s5622,s5623,s5624,s5625,s5626,s5627,s5628,s5629,s5630,s5631,s5632,s5633,s5634,s5635,s5636,s5637,s5638,s5639,s5640,s5641,s5642,s5643,s5644,s5645,s5646,s5647,s5648,s5649,s5650,s5651,s5652,s5653,s5654,s5655,s5656,s5657,s5658,s5659,s5660,s5661,s5662,s5663,s5664,s5665,s5666,s5667,s5668,s5669,s5670,s5671,s5672,s5673,s5674,s5675,s5676,s5677,s5678,s5679,

s5680,s5681,s5682,s5683,s5684,s5685,s5686,s5687,s5688,s5689,s5690,s5691,s5692,s5693,s5694,s5695,s5696,s5697,s5698,s5699,s5700,s5701,s5702,s5703,s5704,s5705,s5706,s5707,s5708,s5709,s5710,s5711,s5712,s5713,s5714,s5715,s5716,s5717,s5718,s5719,s5720,s5721,s5722,s5723,s5724,s5725,s5726,s5727,s5728,s5729,s5730,s5731,s5732,s5733,s5734,s5735,s5736,s5737,s5738,s5739,s5740,s5741,s5742,s5743,s5744,s5745,s5746,s5747,s5748,s5749,s5750,s5751,s5752,s5753,s5754,s5755,s5756,s5757,s5758,s5759,

s5760,s5761,s5762,s5763,s5764,s5765,s5766,s5767,s5768,s5769,s5770,s5771,s5772,s5773,s5774,s5775,s5776,s5777,s5778,s5779,s5780,s5781,s5782,s5783,s5784,s5785,s5786,s5787,s5788,s5789,s5790,s5791,s5792,s5793,s5794,s5795,s5796,s5797,s5798,s5799,s5800,s5801,s5802,s5803,s5804,s5805,s5806,s5807,s5808,s5809,s5810,s5811,s5812,s5813,s5814,s5815,s5816,s5817,s5818,s5819,s5820,s5821,s5822,s5823,s5824,s5825,s5826,s5827,s5828,s5829,s5830,s5831,s5832,s5833,s5834,s5835,s5836,s5837,s5838,s5839,

s5840,s5841,s5842,s5843,s5844,s5845,s5846,s5847,s5848,s5849,s5850,s5851,s5852,s5853,s5854,s5855,s5856,s5857,s5858,s5859,s5860,s5861,s5862,s5863,s5864,s5865,s5866,s5867,s5868,s5869,s5870,s5871,s5872,s5873,s5874,s5875,s5876,s5877,s5878,s5879,s5880,s5881,s5882,s5883,s5884,s5885,s5886,s5887,s5888,s5889,s5890,s5891,s5892,s5893,s5894,s5895,s5896,s5897,s5898,s5899,s5900,s5901,s5902,s5903,s5904,s5905,s5906,s5907,s5908,s5909,s5910,s5911,s5912,s5913,s5914,s5915,s5916,s5917,s5918,s5919,

s5920,s5921,s5922,s5923,s5924,s5925,s5926,s5927,s5928,s5929,s5930,s5931,s5932,s5933,s5934,s5935,s5936,s5937,s5938,s5939,s5940,s5941,s5942,s5943,s5944,s5945,s5946,s5947,s5948,s5949,s5950,s5951,s5952,s5953,s5954,s5955,s5956,s5957,s5958,s5959,s5960,s5961,s5962,s5963,s5964,s5965,s5966,s5967,s5968,s5969,s5970,s5971,s5972,s5973,s5974,s5975,s5976,s5977,s5978,s5979,s5980,s5981,s5982,s5983,s5984,s5985,s5986,s5987,s5988,s5989,s5990,s5991,s5992,s5993,s5994,s5995,s5996,s5997,s5998,s5999,

s6000,s6001,s6002,s6003,s6004,s6005,s6006,s6007,s6008,s6009,s6010,s6011,s6012,s6013,s6014,s6015,s6016,s6017,s6018,s6019,s6020,s6021,s6022,s6023,s6024,s6025,s6026,s6027,s6028,s6029,s6030,s6031,s6032,s6033,s6034,s6035,s6036,s6037,s6038,s6039,s6040,s6041,s6042,s6043,s6044,s6045,s6046,s6047,s6048,s6049,s6050,s6051,s6052,s6053,s6054,s6055,s6056,s6057,s6058,s6059,s6060,s6061,s6062,s6063,s6064,s6065,s6066,s6067,s6068,s6069,s6070,s6071,s6072,s6073,s6074,s6075,s6076,s6077,s6078,s6079,

s6080,s6081,s6082,s6083,s6084,s6085,s6086,s6087,s6088,s6089,s6090,s6091,s6092,s6093,s6094,s6095,s6096,s6097,s6098,s6099,s6100,s6101,s6102,s6103,s6104,s6105,s6106,s6107,s6108,s6109,s6110,s6111,s6112,s6113,s6114,s6115,s6116,s6117,s6118,s6119,s6120,s6121,s6122,s6123,s6124,s6125,s6126,s6127,s6128,s6129,s6130,s6131,s6132,s6133,s6134,s6135,s6136,s6137,s6138,s6139,s6140,s6141,s6142,s6143,s6144,s6145,s6146,s6147,s6148,s6149,s6150,s6151,s6152,s6153,s6154,s6155,s6156,s6157,s6158,s6159,

s6160,s6161,s6162,s6163,s6164,s6165,s6166,s6167,s6168,s6169,s6170,s6171,s6172,s6173,s6174,s6175,s6176,s6177,s6178,s6179,s6180,s6181,s6182,s6183,s6184,s6185,s6186,s6187,s6188,s6189,s6190,s6191,s6192,s6193,s6194,s6195,s6196,s6197,s6198,s6199,s6200,s6201,s6202,s6203,s6204,s6205,s6206,s6207,s6208,s6209,s6210,s6211,s6212,s6213,s6214,s6215,s6216,s6217,s6218,s6219,s6220,s6221,s6222,s6223,s6224,s6225,s6226,s6227,s6228,s6229,s6230,s6231,s6232,s6233,s6234,s6235,s6236,s6237,s6238,s6239,

s6240,s6241,s6242,s6243,s6244,s6245,s6246,s6247,s6248,s6249,s6250,s6251,s6252,s6253,s6254,s6255,s6256,s6257,s6258,s6259,s6260,s6261,s6262,s6263,s6264,s6265,s6266,s6267,s6268,s6269,s6270,s6271,s6272,s6273,s6274,s6275,s6276,s6277,s6278,s6279,s6280,s6281,s6282,s6283,s6284,s6285,s6286,s6287,s6288,s6289,s6290,s6291,s6292,s6293,s6294,s6295,s6296,s6297,s6298,s6299,s6300,s6301,s6302,s6303,s6304,s6305,s6306,s6307,s6308,s6309,s6310,s6311,s6312,s6313,s6314,s6315,s6316,s6317,s6318,s6319,

s6320,s6321,s6322,s6323,s6324,s6325,s6326,s6327,s6328,s6329,s6330,s6331,s6332,s6333,s6334,s6335,s6336,s6337,s6338,s6339,s6340,s6341,s6342,s6343,s6344,s6345,s6346,s6347,s6348,s6349,s6350,s6351,s6352,s6353,s6354,s6355,s6356,s6357,s6358,s6359,s6360,s6361,s6362,s6363,s6364,s6365,s6366,s6367,s6368,s6369,s6370,s6371,s6372,s6373,s6374,s6375,s6376,s6377,s6378,s6379,s6380,s6381,s6382,s6383,s6384,s6385,s6386,s6387,s6388,s6389,s6390,s6391,s6392,s6393,s6394,s6395,s6396,s6397,s6398,s6399,

s6400,s6401,s6402,s6403,s6404,s6405,s6406,s6407,s6408,s6409,s6410,s6411,s6412,s6413,s6414,s6415,s6416,s6417,s6418,s6419,s6420,s6421,s6422,s6423,s6424,s6425,s6426,s6427,s6428,s6429,s6430,s6431,s6432,s6433,s6434,s6435,s6436,s6437,s6438,s6439,s6440,s6441,s6442,s6443,s6444,s6445,s6446,s6447,s6448,s6449,s6450,s6451,s6452,s6453,s6454,s6455,s6456,s6457,s6458,s6459,s6460,s6461,s6462,s6463,s6464,s6465,s6466,s6467,s6468,s6469,s6470,s6471,s6472,s6473,s6474,s6475,s6476,s6477,s6478,s6479,

s6480,s6481,s6482,s6483,s6484,s6485,s6486,s6487,s6488,s6489,s6490,s6491,s6492,s6493,s6494,s6495,s6496,s6497,s6498,s6499,s6500,s6501,s6502,s6503,s6504,s6505,s6506,s6507,s6508,s6509,s6510,s6511,s6512,s6513,s6514,s6515,s6516,s6517,s6518,s6519,s6520,s6521,s6522,s6523,s6524,s6525,s6526,s6527,s6528,s6529,s6530,s6531,s6532,s6533,s6534,s6535,s6536,s6537,s6538,s6539,s6540,s6541,s6542,s6543,s6544,s6545,s6546,s6547,s6548,s6549,s6550,s6551,s6552,s6553,s6554,s6555,s6556,s6557,s6558,s6559,

s6560,s6561,s6562,s6563,s6564,s6565,s6566,s6567,s6568,s6569,s6570,s6571,s6572,s6573,s6574,s6575,s6576,s6577,s6578,s6579,s6580,s6581,s6582,s6583,s6584,s6585,s6586,s6587,s6588,s6589,s6590,s6591,s6592,s6593,s6594,s6595,s6596,s6597,s6598,s6599,s6600,s6601,s6602,s6603,s6604,s6605,s6606,s6607,s6608,s6609,s6610,s6611,s6612,s6613,s6614,s6615,s6616,s6617,s6618,s6619,s6620,s6621,s6622,s6623,s6624,s6625,s6626,s6627,s6628,s6629,s6630,s6631,s6632,s6633,s6634,s6635,s6636,s6637,s6638,s6639,

s6640,s6641,s6642,s6643,s6644,s6645,s6646,s6647,s6648,s6649,s6650,s6651,s6652,s6653,s6654,s6655,s6656,s6657,s6658,s6659,s6660,s6661,s6662,s6663,s6664,s6665,s6666,s6667,s6668,s6669,s6670,s6671,s6672,s6673,s6674,s6675,s6676,s6677,s6678,s6679,s6680,s6681,s6682,s6683,s6684,s6685,s6686,s6687,s6688,s6689,s6690,s6691,s6692,s6693,s6694,s6695,s6696,s6697,s6698,s6699,s6700,s6701,s6702,s6703,s6704,s6705,s6706,s6707,s6708,s6709,s6710,s6711,s6712,s6713,s6714,s6715,s6716,s6717,s6718,s6719,

s6720,s6721,s6722,s6723,s6724,s6725,s6726,s6727,s6728,s6729,s6730,s6731,s6732,s6733,s6734,s6735,s6736,s6737,s6738,s6739,s6740,s6741,s6742,s6743,s6744,s6745,s6746,s6747,s6748,s6749,s6750,s6751,s6752,s6753,s6754,s6755,s6756,s6757,s6758,s6759,s6760,s6761,s6762,s6763,s6764,s6765,s6766,s6767,s6768,s6769,s6770,s6771,s6772,s6773,s6774,s6775,s6776,s6777,s6778,s6779,s6780,s6781,s6782,s6783,s6784,s6785,s6786,s6787,s6788,s6789,s6790,s6791,s6792,s6793,s6794,s6795,s6796,s6797,s6798,s6799,

s6800,s6801,s6802,s6803,s6804,s6805,s6806,s6807,s6808,s6809,s6810,s6811,s6812,s6813,s6814,s6815,s6816,s6817,s6818,s6819,s6820,s6821,s6822,s6823,s6824,s6825,s6826,s6827,s6828,s6829,s6830,s6831,s6832,s6833,s6834,s6835,s6836,s6837,s6838,s6839,s6840,s6841,s6842,s6843,s6844,s6845,s6846,s6847,s6848,s6849,s6850,s6851,s6852,s6853,s6854,s6855,s6856,s6857,s6858,s6859,s6860,s6861,s6862,s6863,s6864,s6865,s6866,s6867,s6868,s6869,s6870,s6871,s6872,s6873,s6874,s6875,s6876,s6877,s6878,s6879,

s6880,s6881,s6882,s6883,s6884,s6885,s6886,s6887,s6888,s6889,s6890,s6891,s6892,s6893,s6894,s6895,s6896,s6897,s6898,s6899,s6900,s6901,s6902,s6903,s6904,s6905,s6906,s6907,s6908,s6909,s6910,s6911,s6912,s6913,s6914,s6915,s6916,s6917,s6918,s6919,s6920,s6921,s6922,s6923,s6924,s6925,s6926,s6927,s6928,s6929,s6930,s6931,s6932,s6933,s6934,s6935,s6936,s6937,s6938,s6939,s6940,s6941,s6942,s6943,s6944,s6945,s6946,s6947,s6948,s6949,s6950,s6951,s6952,s6953,s6954,s6955,s6956,s6957,s6958,s6959,

s6960,s6961,s6962,s6963,s6964,s6965,s6966,s6967,s6968,s6969,s6970,s6971,s6972,s6973,s6974,s6975,s6976,s6977,s6978,s6979,s6980,s6981,s6982,s6983,s6984,s6985,s6986,s6987,s6988,s6989,s6990,s6991,s6992,s6993,s6994,s6995,s6996,s6997,s6998,s6999,s7000,s7001,s7002,s7003,s7004,s7005,s7006,s7007,s7008,s7009,s7010,s7011,s7012,s7013,s7014,s7015,s7016,s7017,s7018,s7019,s7020,s7021,s7022,s7023,s7024,s7025,s7026,s7027,s7028,s7029,s7030,s7031,s7032,s7033,s7034,s7035,s7036,s7037,s7038,s7039,

s7040,s7041,s7042,s7043,s7044,s7045,s7046,s7047,s7048,s7049,s7050,s7051,s7052,s7053,s7054,s7055,s7056,s7057,s7058,s7059,s7060,s7061,s7062,s7063,s7064,s7065,s7066,s7067,s7068,s7069,s7070,s7071,s7072,s7073,s7074,s7075,s7076,s7077,s7078,s7079,s7080,s7081,s7082,s7083,s7084,s7085,s7086,s7087,s7088,s7089,s7090,s7091,s7092,s7093,s7094,s7095,s7096,s7097,s7098,s7099,s7100,s7101,s7102,s7103,s7104,s7105,s7106,s7107,s7108,s7109,s7110,s7111,s7112,s7113,s7114,s7115,s7116,s7117,s7118,s7119,

s7120,s7121,s7122,s7123,s7124,s7125,s7126,s7127,s7128,s7129,s7130,s7131,s7132,s7133,s7134,s7135,s7136,s7137,s7138,s7139,s7140,s7141,s7142,s7143,s7144,s7145,s7146,s7147,s7148,s7149,s7150,s7151,s7152,s7153,s7154,s7155,s7156,s7157,s7158,s7159,s7160,s7161,s7162,s7163,s7164,s7165,s7166,s7167,s7168,s7169,s7170,s7171,s7172,s7173,s7174,s7175,s7176,s7177,s7178,s7179,s7180,s7181,s7182,s7183,s7184,s7185,s7186,s7187,s7188,s7189,s7190,s7191,s7192,s7193,s7194,s7195,s7196,s7197,s7198,s7199,

s7200,s7201,s7202,s7203,s7204,s7205,s7206,s7207,s7208,s7209,s7210,s7211,s7212,s7213,s7214,s7215,s7216,s7217,s7218,s7219,s7220,s7221,s7222,s7223,s7224,s7225,s7226,s7227,s7228,s7229,s7230,s7231,s7232,s7233,s7234,s7235,s7236,s7237,s7238,s7239,s7240,s7241,s7242,s7243,s7244,s7245,s7246,s7247,s7248,s7249,s7250,s7251,s7252,s7253,s7254,s7255,s7256,s7257,s7258,s7259,s7260,s7261,s7262,s7263,s7264,s7265,s7266,s7267,s7268,s7269,s7270,s7271,s7272,s7273,s7274,s7275,s7276,s7277,s7278,s7279,

s7280,s7281,s7282,s7283,s7284,s7285,s7286,s7287,s7288,s7289,s7290,s7291,s7292,s7293,s7294,s7295,s7296,s7297,s7298,s7299,s7300,s7301,s7302,s7303,s7304,s7305,s7306,s7307,s7308,s7309,s7310,s7311,s7312,s7313,s7314,s7315,s7316,s7317,s7318,s7319,s7320,s7321,s7322,s7323,s7324,s7325,s7326,s7327,s7328,s7329,s7330,s7331,s7332,s7333,s7334,s7335,s7336,s7337,s7338,s7339,s7340,s7341,s7342,s7343,s7344,s7345,s7346,s7347,s7348,s7349,s7350,s7351,s7352,s7353,s7354,s7355,s7356,s7357,s7358,s7359,

s7360,s7361,s7362,s7363,s7364,s7365,s7366,s7367,s7368,s7369,s7370,s7371,s7372,s7373,s7374,s7375,s7376,s7377,s7378,s7379,s7380,s7381,s7382,s7383,s7384,s7385,s7386,s7387,s7388,s7389,s7390,s7391,s7392,s7393,s7394,s7395,s7396,s7397,s7398,s7399,s7400,s7401,s7402,s7403,s7404,s7405,s7406,s7407,s7408,s7409,s7410,s7411,s7412,s7413,s7414,s7415,s7416,s7417,s7418,s7419,s7420,s7421,s7422,s7423,s7424,s7425,s7426,s7427,s7428,s7429,s7430,s7431,s7432,s7433,s7434,s7435,s7436,s7437,s7438,s7439,

s7440,s7441,s7442,s7443,s7444,s7445,s7446,s7447,s7448,s7449,s7450,s7451,s7452,s7453,s7454,s7455,s7456,s7457,s7458,s7459,s7460,s7461,s7462,s7463,s7464,s7465,s7466,s7467,s7468,s7469,s7470,s7471,s7472,s7473,s7474,s7475,s7476,s7477,s7478,s7479,s7480,s7481,s7482,s7483,s7484,s7485,s7486,s7487,s7488,s7489,s7490,s7491,s7492,s7493,s7494,s7495,s7496,s7497,s7498,s7499,s7500,s7501,s7502,s7503,s7504,s7505,s7506,s7507,s7508,s7509,s7510,s7511,s7512,s7513,s7514,s7515,s7516,s7517,s7518,s7519,

s7520,s7521,s7522,s7523,s7524,s7525,s7526,s7527,s7528,s7529,s7530,s7531,s7532,s7533,s7534,s7535,s7536,s7537,s7538,s7539,s7540,s7541,s7542,s7543,s7544,s7545,s7546,s7547,s7548,s7549,s7550,s7551,s7552,s7553,s7554,s7555,s7556,s7557,s7558,s7559,s7560,s7561,s7562,s7563,s7564,s7565,s7566,s7567,s7568,s7569,s7570,s7571,s7572,s7573,s7574,s7575,s7576,s7577,s7578,s7579,s7580,s7581,s7582,s7583,s7584,s7585,s7586,s7587,s7588,s7589,s7590,s7591,s7592,s7593,s7594,s7595,s7596,s7597,s7598,s7599,

s7600,s7601,s7602,s7603,s7604,s7605,s7606,s7607,s7608,s7609,s7610,s7611,s7612,s7613,s7614,s7615,s7616,s7617,s7618,s7619,s7620,s7621,s7622,s7623,s7624,s7625,s7626,s7627,s7628,s7629,s7630,s7631,s7632,s7633,s7634,s7635,s7636,s7637,s7638,s7639,s7640,s7641,s7642,s7643,s7644,s7645,s7646,s7647,s7648,s7649,s7650,s7651,s7652,s7653,s7654,s7655,s7656,s7657,s7658,s7659,s7660,s7661,s7662,s7663,s7664,s7665,s7666,s7667,s7668,s7669,s7670,s7671,s7672,s7673,s7674,s7675,s7676,s7677,s7678,s7679,

s7680,s7681,s7682,s7683,s7684,s7685,s7686,s7687,s7688,s7689,s7690,s7691,s7692,s7693,s7694,s7695,s7696,s7697,s7698,s7699,s7700,s7701,s7702,s7703,s7704,s7705,s7706,s7707,s7708,s7709,s7710,s7711,s7712,s7713,s7714,s7715,s7716,s7717,s7718,s7719,s7720,s7721,s7722,s7723,s7724,s7725,s7726,s7727,s7728,s7729,s7730,s7731,s7732,s7733,s7734,s7735,s7736,s7737,s7738,s7739,s7740,s7741,s7742,s7743,s7744,s7745,s7746,s7747,s7748,s7749,s7750,s7751,s7752,s7753,s7754,s7755,s7756,s7757,s7758,s7759,

s7760,s7761,s7762,s7763,s7764,s7765,s7766,s7767,s7768,s7769,s7770,s7771,s7772,s7773,s7774,s7775,s7776,s7777,s7778,s7779,s7780,s7781,s7782,s7783,s7784,s7785,s7786,s7787,s7788,s7789,s7790,s7791,s7792,s7793,s7794,s7795,s7796,s7797,s7798,s7799,s7800,s7801,s7802,s7803,s7804,s7805,s7806,s7807,s7808,s7809,s7810,s7811,s7812,s7813,s7814,s7815,s7816,s7817,s7818,s7819,s7820,s7821,s7822,s7823,s7824,s7825,s7826,s7827,s7828,s7829,s7830,s7831,s7832,s7833,s7834,s7835,s7836,s7837,s7838,s7839,

s7840,s7841,s7842,s7843,s7844,s7845,s7846,s7847,s7848,s7849,s7850,s7851,s7852,s7853,s7854,s7855,s7856,s7857,s7858,s7859,s7860,s7861,s7862,s7863,s7864,s7865,s7866,s7867,s7868,s7869,s7870,s7871,s7872,s7873,s7874,s7875,s7876,s7877,s7878,s7879,s7880,s7881,s7882,s7883,s7884,s7885,s7886,s7887,s7888,s7889,s7890,s7891,s7892,s7893,s7894,s7895,s7896,s7897,s7898,s7899,s7900,s7901,s7902,s7903,s7904,s7905,s7906,s7907,s7908,s7909,s7910,s7911,s7912,s7913,s7914,s7915,s7916,s7917,s7918,s7919,

s7920,s7921,s7922,s7923,s7924,s7925,s7926,s7927,s7928,s7929,s7930,s7931,s7932,s7933,s7934,s7935,s7936,s7937,s7938,s7939,s7940,s7941,s7942,s7943,s7944,s7945,s7946,s7947,s7948,s7949,s7950,s7951,s7952,s7953,s7954,s7955,s7956,s7957,s7958,s7959,s7960,s7961,s7962,s7963,s7964,s7965,s7966,s7967,s7968,s7969,s7970,s7971,s7972,s7973,s7974,s7975,s7976,s7977,s7978,s7979,s7980,s7981,s7982,s7983,s7984,s7985,s7986,s7987,s7988,s7989,s7990,s7991,s7992,s7993,s7994,s7995,s7996,s7997,s7998,s7999,

s8000,s8001,s8002,s8003,s8004,s8005,s8006,s8007,s8008,s8009,s8010,s8011,s8012,s8013,s8014,s8015,s8016,s8017,s8018,s8019,s8020,s8021,s8022,s8023,s8024,s8025,s8026,s8027,s8028,s8029,s8030,s8031,s8032,s8033,s8034,s8035,s8036,s8037,s8038,s8039,s8040,s8041,s8042,s8043,s8044,s8045,s8046,s8047,s8048,s8049,s8050,s8051,s8052,s8053,s8054,s8055,s8056,s8057,s8058,s8059,s8060,s8061,s8062,s8063,s8064,s8065,s8066,s8067,s8068,s8069,s8070,s8071,s8072,s8073,s8074,s8075,s8076,s8077,s8078,s8079,

s8080,s8081,s8082,s8083,s8084,s8085,s8086,s8087,s8088,s8089,s8090,s8091,s8092,s8093,s8094,s8095,s8096,s8097,s8098,s8099,s8100,s8101,s8102,s8103,s8104,s8105,s8106,s8107,s8108,s8109,s8110,s8111,s8112,s8113,s8114,s8115,s8116,s8117,s8118,s8119,s8120,s8121,s8122,s8123,s8124,s8125,s8126,s8127,s8128,s8129,s8130,s8131,s8132,s8133,s8134,s8135,s8136,s8137,s8138,s8139,s8140,s8141,s8142,s8143,s8144,s8145,s8146,s8147,s8148,s8149,s8150,s8151,s8152,s8153,s8154,s8155,s8156,s8157,s8158,s8159,

s8160,s8161,s8162,s8163,s8164,s8165,s8166,s8167,s8168,s8169,s8170,s8171,s8172,s8173,s8174,s8175,s8176,s8177,s8178,s8179,s8180,s8181,s8182,s8183,s8184,s8185,s8186,s8187,s8188,s8189,s8190,s8191,s8192,s8193,s8194,s8195,s8196,s8197,s8198,s8199,s8200,s8201,s8202,s8203,s8204,s8205,s8206,s8207,s8208,s8209,s8210,s8211,s8212,s8213,s8214,s8215,s8216,s8217,s8218,s8219,s8220,s8221,s8222,s8223,s8224,s8225,s8226,s8227,s8228,s8229,s8230,s8231,s8232,s8233,s8234,s8235,s8236,s8237,s8238,s8239,

s8240,s8241,s8242,s8243,s8244,s8245,s8246,s8247,s8248,s8249,s8250,s8251,s8252,s8253,s8254,s8255,s8256,s8257,s8258,s8259,s8260,s8261,s8262,s8263,s8264,s8265,s8266,s8267,s8268,s8269,s8270,s8271,s8272,s8273,s8274,s8275,s8276,s8277,s8278,s8279,s8280,s8281,s8282,s8283,s8284,s8285,s8286,s8287,s8288,s8289,s8290,s8291,s8292,s8293,s8294,s8295,s8296,s8297,s8298,s8299,s8300,s8301,s8302,s8303,s8304,s8305,s8306,s8307,s8308,s8309,s8310,s8311,s8312,s8313,s8314,s8315,s8316,s8317,s8318,s8319,

s8320,s8321,s8322,s8323,s8324,s8325,s8326,s8327,s8328,s8329,s8330,s8331,s8332,s8333,s8334,s8335,s8336,s8337,s8338,s8339,s8340,s8341,s8342,s8343,s8344,s8345,s8346,s8347,s8348,s8349,s8350,s8351,s8352,s8353,s8354,s8355,s8356,s8357,s8358,s8359,s8360,s8361,s8362,s8363,s8364,s8365,s8366,s8367,s8368,s8369,s8370,s8371,s8372,s8373,s8374,s8375,s8376,s8377,s8378,s8379,s8380,s8381,s8382,s8383,s8384,s8385,s8386,s8387,s8388,s8389,s8390,s8391,s8392,s8393,s8394,s8395,s8396,s8397,s8398,s8399,

s8400,s8401,s8402,s8403,s8404,s8405,s8406,s8407,s8408,s8409,s8410,s8411,s8412,s8413,s8414,s8415,s8416,s8417,s8418,s8419,s8420,s8421,s8422,s8423,s8424,s8425,s8426,s8427,s8428,s8429,s8430,s8431,s8432,s8433,s8434,s8435,s8436,s8437,s8438,s8439,s8440,s8441,s8442,s8443,s8444,s8445,s8446,s8447,s8448,s8449,s8450,s8451,s8452,s8453,s8454,s8455,s8456,s8457,s8458,s8459,s8460,s8461,s8462,s8463,s8464,s8465,s8466,s8467,s8468,s8469,s8470,s8471,s8472,s8473,s8474,s8475,s8476,s8477,s8478,s8479,

s8480,s8481,s8482,s8483,s8484,s8485,s8486,s8487,s8488,s8489,s8490,s8491,s8492,s8493,s8494,s8495,s8496,s8497,s8498,s8499,s8500,s8501,s8502,s8503,s8504,s8505,s8506,s8507,s8508,s8509,s8510,s8511,s8512,s8513,s8514,s8515,s8516,s8517,s8518,s8519,s8520,s8521,s8522,s8523,s8524,s8525,s8526,s8527,s8528,s8529,s8530,s8531,s8532,s8533,s8534,s8535,s8536,s8537,s8538,s8539,s8540,s8541,s8542,s8543,s8544,s8545,s8546,s8547,s8548,s8549,s8550,s8551,s8552,s8553,s8554,s8555,s8556,s8557,s8558,s8559,

s8560,s8561,s8562,s8563,s8564,s8565,s8566,s8567,s8568,s8569,s8570,s8571,s8572,s8573,s8574,s8575,s8576,s8577,s8578,s8579,s8580,s8581,s8582,s8583,s8584,s8585,s8586,s8587,s8588,s8589,s8590,s8591,s8592,s8593,s8594,s8595,s8596,s8597,s8598,s8599,s8600,s8601,s8602,s8603,s8604,s8605,s8606,s8607,s8608,s8609,s8610,s8611,s8612,s8613,s8614,s8615,s8616,s8617,s8618,s8619,s8620,s8621,s8622,s8623,s8624,s8625,s8626,s8627,s8628,s8629,s8630,s8631,s8632,s8633,s8634,s8635,s8636,s8637,s8638,s8639,

s8640,s8641,s8642,s8643,s8644,s8645,s8646,s8647,s8648,s8649,s8650,s8651,s8652,s8653,s8654,s8655,s8656,s8657,s8658,s8659,s8660,s8661,s8662,s8663,s8664,s8665,s8666,s8667,s8668,s8669,s8670,s8671,s8672,s8673,s8674,s8675,s8676,s8677,s8678,s8679,s8680,s8681,s8682,s8683,s8684,s8685,s8686,s8687,s8688,s8689,s8690,s8691,s8692,s8693,s8694,s8695,s8696,s8697,s8698,s8699,s8700,s8701,s8702,s8703,s8704,s8705,s8706,s8707,s8708,s8709,s8710,s8711,s8712,s8713,s8714,s8715,s8716,s8717,s8718,s8719,

s8720,s8721,s8722,s8723,s8724,s8725,s8726,s8727,s8728,s8729,s8730,s8731,s8732,s8733,s8734,s8735,s8736,s8737,s8738,s8739,s8740,s8741,s8742,s8743,s8744,s8745,s8746,s8747,s8748,s8749,s8750,s8751,s8752,s8753,s8754,s8755,s8756,s8757,s8758,s8759,s8760,s8761,s8762,s8763,s8764,s8765,s8766,s8767,s8768,s8769,s8770,s8771,s8772,s8773,s8774,s8775,s8776,s8777,s8778,s8779,s8780,s8781,s8782,s8783,s8784,s8785,s8786,s8787,s8788,s8789,s8790,s8791,s8792,s8793,s8794,s8795,s8796,s8797,s8798,s8799,

s8800,s8801,s8802,s8803,s8804,s8805,s8806,s8807,s8808,s8809,s8810,s8811,s8812,s8813,s8814,s8815,s8816,s8817,s8818,s8819,s8820,s8821,s8822,s8823,s8824,s8825,s8826,s8827,s8828,s8829,s8830,s8831,s8832,s8833,s8834,s8835,s8836,s8837,s8838,s8839,s8840,s8841,s8842,s8843,s8844,s8845,s8846,s8847,s8848,s8849,s8850,s8851,s8852,s8853,s8854,s8855,s8856,s8857,s8858,s8859,s8860,s8861,s8862,s8863,s8864,s8865,s8866,s8867,s8868,s8869,s8870,s8871,s8872,s8873,s8874,s8875,s8876,s8877,s8878,s8879,

s8880,s8881,s8882,s8883,s8884,s8885,s8886,s8887,s8888,s8889,s8890,s8891,s8892,s8893,s8894,s8895,s8896,s8897,s8898,s8899,s8900,s8901,s8902,s8903,s8904,s8905,s8906,s8907,s8908,s8909,s8910,s8911,s8912,s8913,s8914,s8915,s8916,s8917,s8918,s8919,s8920,s8921,s8922,s8923,s8924,s8925,s8926,s8927,s8928,s8929,s8930,s8931,s8932,s8933,s8934,s8935,s8936,s8937,s8938,s8939,s8940,s8941,s8942,s8943,s8944,s8945,s8946,s8947,s8948,s8949,s8950,s8951,s8952,s8953,s8954,s8955,s8956,s8957,s8958,s8959,

s8960,s8961,s8962,s8963,s8964,s8965,s8966,s8967,s8968,s8969,s8970,s8971,s8972,s8973,s8974,s8975,s8976,s8977,s8978,s8979,s8980,s8981,s8982,s8983,s8984,s8985,s8986,s8987,s8988,s8989,s8990,s8991,s8992,s8993,s8994,s8995,s8996,s8997,s8998,s8999,s9000,s9001,s9002,s9003,s9004,s9005,s9006,s9007,s9008,s9009,s9010,s9011,s9012,s9013,s9014,s9015,s9016,s9017,s9018,s9019,s9020,s9021,s9022,s9023,s9024,s9025,s9026,s9027,s9028,s9029,s9030,s9031,s9032,s9033,s9034,s9035,s9036,s9037,s9038,s9039,

s9040,s9041,s9042,s9043,s9044,s9045,s9046,s9047,s9048,s9049,s9050,s9051,s9052,s9053,s9054,s9055,s9056,s9057,s9058,s9059,s9060,s9061,s9062,s9063,s9064,s9065,s9066,s9067,s9068,s9069,s9070,s9071,s9072,s9073,s9074,s9075,s9076,s9077,s9078,s9079,s9080,s9081,s9082,s9083,s9084,s9085,s9086,s9087,s9088,s9089,s9090,s9091,s9092,s9093,s9094,s9095,s9096,s9097,s9098,s9099,s9100,s9101,s9102,s9103,s9104,s9105,s9106,s9107,s9108,s9109,s9110,s9111,s9112,s9113,s9114,s9115,s9116,s9117,s9118,s9119,

s9120,s9121,s9122,s9123,s9124,s9125,s9126,s9127,s9128,s9129,s9130,s9131,s9132,s9133,s9134,s9135,s9136,s9137,s9138,s9139,s9140,s9141,s9142,s9143,s9144,s9145,s9146,s9147,s9148,s9149,s9150,s9151,s9152,s9153,s9154,s9155,s9156,s9157,s9158,s9159,s9160,s9161,s9162,s9163,s9164,s9165,s9166,s9167,s9168,s9169,s9170,s9171,s9172,s9173,s9174,s9175,s9176,s9177,s9178,s9179,s9180,s9181,s9182,s9183,s9184,s9185,s9186,s9187,s9188,s9189,s9190,s9191,s9192,s9193,s9194,s9195,s9196,s9197,s9198,s9199,

s9200,s9201,s9202,s9203,s9204,s9205,s9206,s9207,s9208,s9209,s9210,s9211,s9212,s9213,s9214,s9215,s9216,s9217,s9218,s9219,s9220,s9221,s9222,s9223,s9224,s9225,s9226,s9227,s9228,s9229,s9230,s9231,s9232,s9233,s9234,s9235,s9236,s9237,s9238,s9239,s9240,s9241,s9242,s9243,s9244,s9245,s9246,s9247,s9248,s9249,s9250,s9251,s9252,s9253,s9254,s9255,s9256,s9257,s9258,s9259,s9260,s9261,s9262,s9263,s9264,s9265,s9266,s9267,s9268,s9269,s9270,s9271,s9272,s9273,s9274,s9275,s9276,s9277,s9278,s9279,

s9280,s9281,s9282,s9283,s9284,s9285,s9286,s9287,s9288,s9289,s9290,s9291,s9292,s9293,s9294,s9295,s9296,s9297,s9298,s9299,s9300,s9301,s9302,s9303,s9304,s9305,s9306,s9307,s9308,s9309,s9310,s9311,s9312,s9313,s9314,s9315,s9316,s9317,s9318,s9319,s9320,s9321,s9322,s9323,s9324,s9325,s9326,s9327,s9328,s9329,s9330,s9331,s9332,s9333,s9334,s9335,s9336,s9337,s9338,s9339,s9340,s9341,s9342,s9343,s9344,s9345,s9346,s9347,s9348,s9349,s9350,s9351,s9352,s9353,s9354,s9355,s9356,s9357,s9358,s9359,

s9360,s9361,s9362,s9363,s9364,s9365,s9366,s9367,s9368,s9369,s9370,s9371,s9372,s9373,s9374,s9375,s9376,s9377,s9378,s9379,s9380,s9381,s9382,s9383,s9384,s9385,s9386,s9387,s9388,s9389,s9390,s9391,s9392,s9393,s9394,s9395,s9396,s9397,s9398,s9399,s9400,s9401,s9402,s9403,s9404,s9405,s9406,s9407,s9408,s9409,s9410,s9411,s9412,s9413,s9414,s9415,s9416,s9417,s9418,s9419,s9420,s9421,s9422,s9423,s9424,s9425,s9426,s9427,s9428,s9429,s9430,s9431,s9432,s9433,s9434,s9435,s9436,s9437,s9438,s9439,

s9440,s9441,s9442,s9443,s9444,s9445,s9446,s9447,s9448,s9449,s9450,s9451,s9452,s9453,s9454,s9455,s9456,s9457,s9458,s9459,s9460,s9461,s9462,s9463,s9464,s9465,s9466,s9467,s9468,s9469,s9470,s9471,s9472,s9473,s9474,s9475,s9476,s9477,s9478,s9479,s9480,s9481,s9482,s9483,s9484,s9485,s9486,s9487,s9488,s9489,s9490,s9491,s9492,s9493,s9494,s9495,s9496,s9497,s9498,s9499,s9500,s9501,s9502,s9503,s9504,s9505,s9506,s9507,s9508,s9509,s9510,s9511,s9512,s9513,s9514,s9515,s9516,s9517,s9518,s9519,

s9520,s9521,s9522,s9523,s9524,s9525,s9526,s9527,s9528,s9529,s9530,s9531,s9532,s9533,s9534,s9535,s9536,s9537,s9538,s9539,s9540,s9541,s9542,s9543,s9544,s9545,s9546,s9547,s9548,s9549,s9550,s9551,s9552,s9553,s9554,s9555,s9556,s9557,s9558,s9559,s9560,s9561,s9562,s9563,s9564,s9565,s9566,s9567,s9568,s9569,s9570,s9571,s9572,s9573,s9574,s9575,s9576,s9577,s9578,s9579,s9580,s9581,s9582,s9583,s9584,s9585,s9586,s9587,s9588,s9589,s9590,s9591,s9592,s9593,s9594,s9595,s9596,s9597,s9598,s9599,

s9600,s9601,s9602,s9603,s9604,s9605,s9606,s9607,s9608,s9609,s9610,s9611,s9612,s9613,s9614,s9615,s9616,s9617,s9618,s9619,s9620,s9621,s9622,s9623,s9624,s9625,s9626,s9627,s9628,s9629,s9630,s9631,s9632,s9633,s9634,s9635,s9636,s9637,s9638,s9639,s9640,s9641,s9642,s9643,s9644,s9645,s9646,s9647,s9648,s9649,s9650,s9651,s9652,s9653,s9654,s9655,s9656,s9657,s9658,s9659,s9660,s9661,s9662,s9663,s9664,s9665,s9666,s9667,s9668,s9669,s9670,s9671,s9672,s9673,s9674,s9675,s9676,s9677,s9678,s9679,

s9680,s9681,s9682,s9683,s9684,s9685,s9686,s9687,s9688,s9689,s9690,s9691,s9692,s9693,s9694,s9695,s9696,s9697,s9698,s9699,s9700,s9701,s9702,s9703,s9704,s9705,s9706,s9707,s9708,s9709,s9710,s9711,s9712,s9713,s9714,s9715,s9716,s9717,s9718,s9719,s9720,s9721,s9722,s9723,s9724,s9725,s9726,s9727,s9728,s9729,s9730,s9731,s9732,s9733,s9734,s9735,s9736,s9737,s9738,s9739,s9740,s9741,s9742,s9743,s9744,s9745,s9746,s9747,s9748,s9749,s9750,s9751,s9752,s9753,s9754,s9755,s9756,s9757,s9758,s9759,

s9760,s9761,s9762,s9763,s9764,s9765,s9766,s9767,s9768,s9769,s9770,s9771,s9772,s9773,s9774,s9775,s9776,s9777,s9778,s9779,s9780,s9781,s9782,s9783,s9784,s9785,s9786,s9787,s9788,s9789,s9790,s9791,s9792,s9793,s9794,s9795,s9796,s9797,s9798,s9799,s9800,s9801,s9802,s9803,s9804,s9805,s9806,s9807,s9808,s9809,s9810,s9811,s9812,s9813,s9814,s9815,s9816,s9817,s9818,s9819,s9820,s9821,s9822,s9823,s9824,s9825,s9826,s9827,s9828,s9829,s9830,s9831,s9832,s9833,s9834,s9835,s9836,s9837,s9838,s9839,

s9840,s9841,s9842,s9843,s9844,s9845,s9846,s9847,s9848,s9849,s9850,s9851,s9852,s9853,s9854,s9855,s9856,s9857,s9858,s9859,s9860,s9861,s9862,s9863,s9864,s9865,s9866,s9867,s9868,s9869,s9870,s9871,s9872,s9873,s9874,s9875,s9876,s9877,s9878,s9879,s9880,s9881,s9882,s9883,s9884,s9885,s9886,s9887,s9888,s9889,s9890,s9891,s9892,s9893,s9894,s9895,s9896,s9897,s9898,s9899,s9900,s9901,s9902,s9903,s9904,s9905,s9906,s9907,s9908,s9909,s9910,s9911,s9912,s9913,s9914,s9915,s9916,s9917,s9918,s9919,

s9920,s9921,s9922,s9923,s9924,s9925,s9926,s9927,s9928,s9929,s9930,s9931,s9932,s9933,s9934,s9935,s9936,s9937,s9938,s9939,s9940,s9941,s9942,s9943,s9944,s9945,s9946,s9947,s9948,s9949,s9950,s9951,s9952,s9953,s9954,s9955,s9956,s9957,s9958,s9959,s9960,s9961,s9962,s9963,s9964,s9965,s9966,s9967,s9968,s9969,s9970,s9971,s9972,s9973,s9974,s9975,s9976,s9977,s9978,s9979,s9980,s9981,s9982,s9983,s9984,s9985,s9986,s9987,s9988,s9989,s9990,s9991,s9992,s9993,s9994,s9995,s9996,s9997,s9998,s9999,

s10000,s10001,s10002,s10003,s10004,s10005,s10006,s10007,s10008,s10009,s10010,s10011,s10012,s10013,s10014,s10015,s10016,s10017,s10018,s10019,s10020,s10021,s10022,s10023,s10024,s10025,s10026,s10027,s10028,s10029,s10030,s10031,s10032,s10033,s10034,s10035,s10036,s10037,s10038,s10039,s10040,s10041,s10042,s10043,s10044,s10045,s10046,s10047,s10048,s10049,s10050,s10051,s10052,s10053,s10054,s10055,s10056,s10057,s10058,s10059,s10060,s10061,s10062,s10063,s10064,s10065,s10066,s10067,s10068,s10069,s10070,s10071,s10072,s10073,s10074,s10075,s10076,s10077,s10078,s10079,

s10080,s10081,s10082,s10083,s10084,s10085,s10086,s10087,s10088,s10089,s10090,s10091,s10092,s10093,s10094,s10095,s10096,s10097,s10098,s10099,s10100,s10101,s10102,s10103,s10104,s10105,s10106,s10107,s10108,s10109,s10110,s10111,s10112,s10113,s10114,s10115,s10116,s10117,s10118,s10119,s10120,s10121,s10122,s10123,s10124,s10125,s10126,s10127,s10128,s10129,s10130,s10131,s10132,s10133,s10134,s10135,s10136,s10137,s10138,s10139,s10140,s10141,s10142,s10143,s10144,s10145,s10146,s10147,s10148,s10149,s10150,s10151,s10152,s10153,s10154,s10155,s10156,s10157,s10158,s10159,

s10160,s10161,s10162,s10163,s10164,s10165,s10166,s10167,s10168,s10169,s10170,s10171,s10172,s10173,s10174,s10175,s10176,s10177,s10178,s10179,s10180,s10181,s10182,s10183,s10184,s10185,s10186,s10187,s10188,s10189,s10190,s10191,s10192,s10193,s10194,s10195,s10196,s10197,s10198,s10199,s10200,s10201,s10202,s10203,s10204,s10205,s10206,s10207,s10208,s10209,s10210,s10211,s10212,s10213,s10214,s10215,s10216,s10217,s10218,s10219,s10220,s10221,s10222,s10223,s10224,s10225,s10226,s10227,s10228,s10229,s10230,s10231,s10232,s10233,s10234,s10235,s10236,s10237,s10238,s10239,

s10240,s10241,s10242,s10243,s10244,s10245,s10246,s10247,s10248,s10249,s10250,s10251,s10252,s10253,s10254,s10255,s10256,s10257,s10258,s10259,s10260,s10261,s10262,s10263,s10264,s10265,s10266,s10267,s10268,s10269,s10270,s10271,s10272,s10273,s10274,s10275,s10276,s10277,s10278,s10279,s10280,s10281,s10282,s10283,s10284,s10285,s10286,s10287,s10288,s10289,s10290,s10291,s10292,s10293,s10294,s10295,s10296,s10297,s10298,s10299,s10300,s10301,s10302,s10303,s10304,s10305,s10306,s10307,s10308,s10309,s10310,s10311,s10312,s10313,s10314,s10315,s10316,s10317,s10318,s10319,

s10320,s10321,s10322,s10323,s10324,s10325,s10326,s10327,s10328,s10329,s10330,s10331,s10332,s10333,s10334,s10335,s10336,s10337,s10338,s10339,s10340,s10341,s10342,s10343,s10344,s10345,s10346,s10347,s10348,s10349,s10350,s10351,s10352,s10353,s10354,s10355,s10356,s10357,s10358,s10359,s10360,s10361,s10362,s10363,s10364,s10365,s10366,s10367,s10368,s10369,s10370,s10371,s10372,s10373,s10374,s10375,s10376,s10377,s10378,s10379,s10380,s10381,s10382,s10383,s10384,s10385,s10386,s10387,s10388,s10389,s10390,s10391,s10392,s10393,s10394,s10395,s10396,s10397,s10398,s10399,

s10400,s10401,s10402,s10403,s10404,s10405,s10406,s10407,s10408,s10409,s10410,s10411,s10412,s10413,s10414,s10415,s10416,s10417,s10418,s10419,s10420,s10421,s10422,s10423,s10424,s10425,s10426,s10427,s10428,s10429,s10430,s10431,s10432,s10433,s10434,s10435,s10436,s10437,s10438,s10439,s10440,s10441,s10442,s10443,s10444,s10445,s10446,s10447,s10448,s10449,s10450,s10451,s10452,s10453,s10454,s10455,s10456,s10457,s10458,s10459,s10460,s10461,s10462,s10463,s10464,s10465,s10466,s10467,s10468,s10469,s10470,s10471,s10472,s10473,s10474,s10475,s10476,s10477,s10478,s10479,

s10480,s10481,s10482,s10483,s10484,s10485,s10486,s10487,s10488,s10489,s10490,s10491,s10492,s10493,s10494,s10495,s10496,s10497,s10498,s10499,s10500,s10501,s10502,s10503,s10504,s10505,s10506,s10507,s10508,s10509,s10510,s10511,s10512,s10513,s10514,s10515,s10516,s10517,s10518,s10519,s10520,s10521,s10522,s10523,s10524,s10525,s10526,s10527,s10528,s10529,s10530,s10531,s10532,s10533,s10534,s10535,s10536,s10537,s10538,s10539,s10540,s10541,s10542,s10543,s10544,s10545,s10546,s10547,s10548,s10549,s10550,s10551,s10552,s10553,s10554,s10555,s10556,s10557,s10558,s10559,

s10560,s10561,s10562,s10563,s10564,s10565,s10566,s10567,s10568,s10569,s10570,s10571,s10572,s10573,s10574,s10575,s10576,s10577,s10578,s10579,s10580,s10581,s10582,s10583,s10584,s10585,s10586,s10587,s10588,s10589,s10590,s10591,s10592,s10593,s10594,s10595,s10596,s10597,s10598,s10599,s10600,s10601,s10602,s10603,s10604,s10605,s10606,s10607,s10608,s10609,s10610,s10611,s10612,s10613,s10614,s10615,s10616,s10617,s10618,s10619,s10620,s10621,s10622,s10623,s10624,s10625,s10626,s10627,s10628,s10629,s10630,s10631,s10632,s10633,s10634,s10635,s10636,s10637,s10638,s10639,

s10640,s10641,s10642,s10643,s10644,s10645,s10646,s10647,s10648,s10649,s10650,s10651,s10652,s10653,s10654,s10655,s10656,s10657,s10658,s10659,s10660,s10661,s10662,s10663,s10664,s10665,s10666,s10667,s10668,s10669,s10670,s10671,s10672,s10673,s10674,s10675,s10676,s10677,s10678,s10679,s10680,s10681,s10682,s10683,s10684,s10685,s10686,s10687,s10688,s10689,s10690,s10691,s10692,s10693,s10694,s10695,s10696,s10697,s10698,s10699,s10700,s10701,s10702,s10703,s10704,s10705,s10706,s10707,s10708,s10709,s10710,s10711,s10712,s10713,s10714,s10715,s10716,s10717,s10718,s10719,

s10720,s10721,s10722,s10723,s10724,s10725,s10726,s10727,s10728,s10729,s10730,s10731,s10732,s10733,s10734,s10735,s10736,s10737,s10738,s10739,s10740,s10741,s10742,s10743,s10744,s10745,s10746,s10747,s10748,s10749,s10750,s10751,s10752,s10753,s10754,s10755,s10756,s10757,s10758,s10759,s10760,s10761,s10762,s10763,s10764,s10765,s10766,s10767,s10768,s10769,s10770,s10771,s10772,s10773,s10774,s10775,s10776,s10777,s10778,s10779,s10780,s10781,s10782,s10783,s10784,s10785,s10786,s10787,s10788,s10789,s10790,s10791,s10792,s10793,s10794,s10795,s10796,s10797,s10798,s10799,

s10800,s10801,s10802,s10803,s10804,s10805,s10806,s10807,s10808,s10809,s10810,s10811,s10812,s10813,s10814,s10815,s10816,s10817,s10818,s10819,s10820,s10821,s10822,s10823,s10824,s10825,s10826,s10827,s10828,s10829,s10830,s10831,s10832,s10833,s10834,s10835,s10836,s10837,s10838,s10839,s10840,s10841,s10842,s10843,s10844,s10845,s10846,s10847,s10848,s10849,s10850,s10851,s10852,s10853,s10854,s10855,s10856,s10857,s10858,s10859,s10860,s10861,s10862,s10863,s10864,s10865,s10866,s10867,s10868,s10869,s10870,s10871,s10872,s10873,s10874,s10875,s10876,s10877,s10878,s10879,

s10880,s10881,s10882,s10883,s10884,s10885,s10886,s10887,s10888,s10889,s10890,s10891,s10892,s10893,s10894,s10895,s10896,s10897,s10898,s10899,s10900,s10901,s10902,s10903,s10904,s10905,s10906,s10907,s10908,s10909,s10910,s10911,s10912,s10913,s10914,s10915,s10916,s10917,s10918,s10919,s10920,s10921,s10922,s10923,s10924,s10925,s10926,s10927,s10928,s10929,s10930,s10931,s10932,s10933,s10934,s10935,s10936,s10937,s10938,s10939,s10940,s10941,s10942,s10943,s10944,s10945,s10946,s10947,s10948,s10949,s10950,s10951,s10952,s10953,s10954,s10955,s10956,s10957,s10958,s10959,

s10960,s10961,s10962,s10963,s10964,s10965,s10966,s10967,s10968,s10969,s10970,s10971,s10972,s10973,s10974,s10975,s10976,s10977,s10978,s10979,s10980,s10981,s10982,s10983,s10984,s10985,s10986,s10987,s10988,s10989,s10990,s10991,s10992,s10993,s10994,s10995,s10996,s10997,s10998,s10999,s11000,s11001,s11002,s11003,s11004,s11005,s11006,s11007,s11008,s11009,s11010,s11011,s11012,s11013,s11014,s11015,s11016,s11017,s11018,s11019,s11020,s11021,s11022,s11023,s11024,s11025,s11026,s11027,s11028,s11029,s11030,s11031,s11032,s11033,s11034,s11035,s11036,s11037,s11038,s11039,

s11040,s11041,s11042,s11043,s11044,s11045,s11046,s11047,s11048,s11049,s11050,s11051,s11052,s11053,s11054,s11055,s11056,s11057,s11058,s11059,s11060,s11061,s11062,s11063,s11064,s11065,s11066,s11067,s11068,s11069,s11070,s11071,s11072,s11073,s11074,s11075,s11076,s11077,s11078,s11079,s11080,s11081,s11082,s11083,s11084,s11085,s11086,s11087,s11088,s11089,s11090,s11091,s11092,s11093,s11094,s11095,s11096,s11097,s11098,s11099,s11100,s11101,s11102,s11103,s11104,s11105,s11106,s11107,s11108,s11109,s11110,s11111,s11112,s11113,s11114,s11115,s11116,s11117,s11118,s11119,

s11120,s11121,s11122,s11123,s11124,s11125,s11126,s11127,s11128,s11129,s11130,s11131,s11132,s11133,s11134,s11135,s11136,s11137,s11138,s11139,s11140,s11141,s11142,s11143,s11144,s11145,s11146,s11147,s11148,s11149,s11150,s11151,s11152,s11153,s11154,s11155,s11156,s11157,s11158,s11159,s11160,s11161,s11162,s11163,s11164,s11165,s11166,s11167,s11168,s11169,s11170,s11171,s11172,s11173,s11174,s11175,s11176,s11177,s11178,s11179,s11180,s11181,s11182,s11183,s11184,s11185,s11186,s11187,s11188,s11189,s11190,s11191,s11192,s11193,s11194,s11195,s11196,s11197,s11198,s11199,

s11200,s11201,s11202,s11203,s11204,s11205,s11206,s11207,s11208,s11209,s11210,s11211,s11212,s11213,s11214,s11215,s11216,s11217,s11218,s11219,s11220,s11221,s11222,s11223,s11224,s11225,s11226,s11227,s11228,s11229,s11230,s11231,s11232,s11233,s11234,s11235,s11236,s11237,s11238,s11239,s11240,s11241,s11242,s11243,s11244,s11245,s11246,s11247,s11248,s11249,s11250,s11251,s11252,s11253,s11254,s11255,s11256,s11257,s11258,s11259,s11260,s11261,s11262,s11263,s11264,s11265,s11266,s11267,s11268,s11269,s11270,s11271,s11272,s11273,s11274,s11275,s11276,s11277,s11278,s11279,

s11280,s11281,s11282,s11283,s11284,s11285,s11286,s11287,s11288,s11289,s11290,s11291,s11292,s11293,s11294,s11295,s11296,s11297,s11298,s11299,s11300,s11301,s11302,s11303,s11304,s11305,s11306,s11307,s11308,s11309,s11310,s11311,s11312,s11313,s11314,s11315,s11316,s11317,s11318,s11319,s11320,s11321,s11322,s11323,s11324,s11325,s11326,s11327,s11328,s11329,s11330,s11331,s11332,s11333,s11334,s11335,s11336,s11337,s11338,s11339,s11340,s11341,s11342,s11343,s11344,s11345,s11346,s11347,s11348,s11349,s11350,s11351,s11352,s11353,s11354,s11355,s11356,s11357,s11358,s11359,

s11360,s11361,s11362,s11363,s11364,s11365,s11366,s11367,s11368,s11369,s11370,s11371,s11372,s11373,s11374,s11375,s11376,s11377,s11378,s11379,s11380,s11381,s11382,s11383,s11384,s11385,s11386,s11387,s11388,s11389,s11390,s11391,s11392,s11393,s11394,s11395,s11396,s11397,s11398,s11399,s11400,s11401,s11402,s11403,s11404,s11405,s11406,s11407,s11408,s11409,s11410,s11411,s11412,s11413,s11414,s11415,s11416,s11417,s11418,s11419,s11420,s11421,s11422,s11423,s11424,s11425,s11426,s11427,s11428,s11429,s11430,s11431,s11432,s11433,s11434,s11435,s11436,s11437,s11438,s11439,

s11440,s11441,s11442,s11443,s11444,s11445,s11446,s11447,s11448,s11449,s11450,s11451,s11452,s11453,s11454,s11455,s11456,s11457,s11458,s11459,s11460,s11461,s11462,s11463,s11464,s11465,s11466,s11467,s11468,s11469,s11470,s11471,s11472,s11473,s11474,s11475,s11476,s11477,s11478,s11479,s11480,s11481,s11482,s11483,s11484,s11485,s11486,s11487,s11488,s11489,s11490,s11491,s11492,s11493,s11494,s11495,s11496,s11497,s11498,s11499,s11500,s11501,s11502,s11503,s11504,s11505,s11506,s11507,s11508,s11509,s11510,s11511,s11512,s11513,s11514,s11515,s11516,s11517,s11518,s11519,

s11520,s11521,s11522,s11523,s11524,s11525,s11526,s11527,s11528,s11529,s11530,s11531,s11532,s11533,s11534,s11535,s11536,s11537,s11538,s11539,s11540,s11541,s11542,s11543,s11544,s11545,s11546,s11547,s11548,s11549,s11550,s11551,s11552,s11553,s11554,s11555,s11556,s11557,s11558,s11559,s11560,s11561,s11562,s11563,s11564,s11565,s11566,s11567,s11568,s11569,s11570,s11571,s11572,s11573,s11574,s11575,s11576,s11577,s11578,s11579,s11580,s11581,s11582,s11583,s11584,s11585,s11586,s11587,s11588,s11589,s11590,s11591,s11592,s11593,s11594,s11595,s11596,s11597,s11598,s11599,

s11600,s11601,s11602,s11603,s11604,s11605,s11606,s11607,s11608,s11609,s11610,s11611,s11612,s11613,s11614,s11615,s11616,s11617,s11618,s11619,s11620,s11621,s11622,s11623,s11624,s11625,s11626,s11627,s11628,s11629,s11630,s11631,s11632,s11633,s11634,s11635,s11636,s11637,s11638,s11639,s11640,s11641,s11642,s11643,s11644,s11645,s11646,s11647,s11648,s11649,s11650,s11651,s11652,s11653,s11654,s11655,s11656,s11657,s11658,s11659,s11660,s11661,s11662,s11663,s11664,s11665,s11666,s11667,s11668,s11669,s11670,s11671,s11672,s11673,s11674,s11675,s11676,s11677,s11678,s11679,

s11680,s11681,s11682,s11683,s11684,s11685,s11686,s11687,s11688,s11689,s11690,s11691,s11692,s11693,s11694,s11695,s11696,s11697,s11698,s11699,s11700,s11701,s11702,s11703,s11704,s11705,s11706,s11707,s11708,s11709,s11710,s11711,s11712,s11713,s11714,s11715,s11716,s11717,s11718,s11719,s11720,s11721,s11722,s11723,s11724,s11725,s11726,s11727,s11728,s11729,s11730,s11731,s11732,s11733,s11734,s11735,s11736,s11737,s11738,s11739,s11740,s11741,s11742,s11743,s11744,s11745,s11746,s11747,s11748,s11749,s11750,s11751,s11752,s11753,s11754,s11755,s11756,s11757,s11758,s11759,

s11760,s11761,s11762,s11763,s11764,s11765,s11766,s11767,s11768,s11769,s11770,s11771,s11772,s11773,s11774,s11775,s11776,s11777,s11778,s11779,s11780,s11781,s11782,s11783,s11784,s11785,s11786,s11787,s11788,s11789,s11790,s11791,s11792,s11793,s11794,s11795,s11796,s11797,s11798,s11799,s11800,s11801,s11802,s11803,s11804,s11805,s11806,s11807,s11808,s11809,s11810,s11811,s11812,s11813,s11814,s11815,s11816,s11817,s11818,s11819,s11820,s11821,s11822,s11823,s11824,s11825,s11826,s11827,s11828,s11829,s11830,s11831,s11832,s11833,s11834,s11835,s11836,s11837,s11838,s11839,

s11840,s11841,s11842,s11843,s11844,s11845,s11846,s11847,s11848,s11849,s11850,s11851,s11852,s11853,s11854,s11855,s11856,s11857,s11858,s11859,s11860,s11861,s11862,s11863,s11864,s11865,s11866,s11867,s11868,s11869,s11870,s11871,s11872,s11873,s11874,s11875,s11876,s11877,s11878,s11879,s11880,s11881,s11882,s11883,s11884,s11885,s11886,s11887,s11888,s11889,s11890,s11891,s11892,s11893,s11894,s11895,s11896,s11897,s11898,s11899,s11900,s11901,s11902,s11903,s11904,s11905,s11906,s11907,s11908,s11909,s11910,s11911,s11912,s11913,s11914,s11915,s11916,s11917,s11918,s11919,

s11920,s11921,s11922,s11923,s11924,s11925,s11926,s11927,s11928,s11929,s11930,s11931,s11932,s11933,s11934,s11935,s11936,s11937,s11938,s11939,s11940,s11941,s11942,s11943,s11944,s11945,s11946,s11947,s11948,s11949,s11950,s11951,s11952,s11953,s11954,s11955,s11956,s11957,s11958,s11959,s11960,s11961,s11962,s11963,s11964,s11965,s11966,s11967,s11968,s11969,s11970,s11971,s11972,s11973,s11974,s11975,s11976,s11977,s11978,s11979,s11980,s11981,s11982,s11983,s11984,s11985,s11986,s11987,s11988,s11989,s11990,s11991,s11992,s11993,s11994,s11995,s11996,s11997,s11998,s11999,

s12000,s12001,s12002,s12003,s12004,s12005,s12006,s12007,s12008,s12009,s12010,s12011,s12012,s12013,s12014,s12015,s12016,s12017,s12018,s12019,s12020,s12021,s12022,s12023,s12024,s12025,s12026,s12027,s12028,s12029,s12030,s12031,s12032,s12033,s12034,s12035,s12036,s12037,s12038,s12039,s12040,s12041,s12042,s12043,s12044,s12045,s12046,s12047,s12048,s12049,s12050,s12051,s12052,s12053,s12054,s12055,s12056,s12057,s12058,s12059,s12060,s12061,s12062,s12063,s12064,s12065,s12066,s12067,s12068,s12069,s12070,s12071,s12072,s12073,s12074,s12075,s12076,s12077,s12078,s12079,

s12080,s12081,s12082,s12083,s12084,s12085,s12086,s12087,s12088,s12089,s12090,s12091,s12092,s12093,s12094,s12095,s12096,s12097,s12098,s12099,s12100,s12101,s12102,s12103,s12104,s12105,s12106,s12107,s12108,s12109,s12110,s12111,s12112,s12113,s12114,s12115,s12116,s12117,s12118,s12119,s12120,s12121,s12122,s12123,s12124,s12125,s12126,s12127,s12128,s12129,s12130,s12131,s12132,s12133,s12134,s12135,s12136,s12137,s12138,s12139,s12140,s12141,s12142,s12143,s12144,s12145,s12146,s12147,s12148,s12149,s12150,s12151,s12152,s12153,s12154,s12155,s12156,s12157,s12158,s12159,

s12160,s12161,s12162,s12163,s12164,s12165,s12166,s12167,s12168,s12169,s12170,s12171,s12172,s12173,s12174,s12175,s12176,s12177,s12178,s12179,s12180,s12181,s12182,s12183,s12184,s12185,s12186,s12187,s12188,s12189,s12190,s12191,s12192,s12193,s12194,s12195,s12196,s12197,s12198,s12199,s12200,s12201,s12202,s12203,s12204,s12205,s12206,s12207,s12208,s12209,s12210,s12211,s12212,s12213,s12214,s12215,s12216,s12217,s12218,s12219,s12220,s12221,s12222,s12223,s12224,s12225,s12226,s12227,s12228,s12229,s12230,s12231,s12232,s12233,s12234,s12235,s12236,s12237,s12238,s12239,

s12240,s12241,s12242,s12243,s12244,s12245,s12246,s12247,s12248,s12249,s12250,s12251,s12252,s12253,s12254,s12255,s12256,s12257,s12258,s12259,s12260,s12261,s12262,s12263,s12264,s12265,s12266,s12267,s12268,s12269,s12270,s12271,s12272,s12273,s12274,s12275,s12276,s12277,s12278,s12279,s12280,s12281,s12282,s12283,s12284,s12285,s12286,s12287,s12288,s12289,s12290,s12291,s12292,s12293,s12294,s12295,s12296,s12297,s12298,s12299,s12300,s12301,s12302,s12303,s12304,s12305,s12306,s12307,s12308,s12309,s12310,s12311,s12312,s12313,s12314,s12315,s12316,s12317,s12318,s12319,

s12320,s12321,s12322,s12323,s12324,s12325,s12326,s12327,s12328,s12329,s12330,s12331,s12332,s12333,s12334,s12335,s12336,s12337,s12338,s12339,s12340,s12341,s12342,s12343,s12344,s12345,s12346,s12347,s12348,s12349,s12350,s12351,s12352,s12353,s12354,s12355,s12356,s12357,s12358,s12359,s12360,s12361,s12362,s12363,s12364,s12365,s12366,s12367,s12368,s12369,s12370,s12371,s12372,s12373,s12374,s12375,s12376,s12377,s12378,s12379,s12380,s12381,s12382,s12383,s12384,s12385,s12386,s12387,s12388,s12389,s12390,s12391,s12392,s12393,s12394,s12395,s12396,s12397,s12398,s12399,

s12400,s12401,s12402,s12403,s12404,s12405,s12406,s12407,s12408,s12409,s12410,s12411,s12412,s12413,s12414,s12415,s12416,s12417,s12418,s12419,s12420,s12421,s12422,s12423,s12424,s12425,s12426,s12427,s12428,s12429,s12430,s12431,s12432,s12433,s12434,s12435,s12436,s12437,s12438,s12439,s12440,s12441,s12442,s12443,s12444,s12445,s12446,s12447,s12448,s12449,s12450,s12451,s12452,s12453,s12454,s12455,s12456,s12457,s12458,s12459,s12460,s12461,s12462,s12463,s12464,s12465,s12466,s12467,s12468,s12469,s12470,s12471,s12472,s12473,s12474,s12475,s12476,s12477,s12478,s12479,

s12480,s12481,s12482,s12483,s12484,s12485,s12486,s12487,s12488,s12489,s12490,s12491,s12492,s12493,s12494,s12495,s12496,s12497,s12498,s12499,s12500,s12501,s12502,s12503,s12504,s12505,s12506,s12507,s12508,s12509,s12510,s12511,s12512,s12513,s12514,s12515,s12516,s12517,s12518,s12519,s12520,s12521,s12522,s12523,s12524,s12525,s12526,s12527,s12528,s12529,s12530,s12531,s12532,s12533,s12534,s12535,s12536,s12537,s12538,s12539,s12540,s12541,s12542,s12543,s12544,s12545,s12546,s12547,s12548,s12549,s12550,s12551,s12552,s12553,s12554,s12555,s12556,s12557,s12558,s12559,

s12560,s12561,s12562,s12563,s12564,s12565,s12566,s12567,s12568,s12569,s12570,s12571,s12572,s12573,s12574,s12575,s12576,s12577,s12578,s12579,s12580,s12581,s12582,s12583,s12584,s12585,s12586,s12587,s12588,s12589,s12590,s12591,s12592,s12593,s12594,s12595,s12596,s12597,s12598,s12599,s12600,s12601,s12602,s12603,s12604,s12605,s12606,s12607,s12608,s12609,s12610,s12611,s12612,s12613,s12614,s12615,s12616,s12617,s12618,s12619,s12620,s12621,s12622,s12623,s12624,s12625,s12626,s12627,s12628,s12629,s12630,s12631,s12632,s12633,s12634,s12635,s12636,s12637,s12638,s12639,

s12640,s12641,s12642,s12643,s12644,s12645,s12646,s12647,s12648,s12649,s12650,s12651,s12652,s12653,s12654,s12655,s12656,s12657,s12658,s12659,s12660,s12661,s12662,s12663,s12664,s12665,s12666,s12667,s12668,s12669,s12670,s12671,s12672,s12673,s12674,s12675,s12676,s12677,s12678,s12679,s12680,s12681,s12682,s12683,s12684,s12685,s12686,s12687,s12688,s12689,s12690,s12691,s12692,s12693,s12694,s12695,s12696,s12697,s12698,s12699,s12700,s12701,s12702,s12703,s12704,s12705,s12706,s12707,s12708,s12709,s12710,s12711,s12712,s12713,s12714,s12715,s12716,s12717,s12718,s12719,

s12720,s12721,s12722,s12723,s12724,s12725,s12726,s12727,s12728,s12729,s12730,s12731,s12732,s12733,s12734,s12735,s12736,s12737,s12738,s12739,s12740,s12741,s12742,s12743,s12744,s12745,s12746,s12747,s12748,s12749,s12750,s12751,s12752,s12753,s12754,s12755,s12756,s12757,s12758,s12759,s12760,s12761,s12762,s12763,s12764,s12765,s12766,s12767,s12768,s12769,s12770,s12771,s12772,s12773,s12774,s12775,s12776,s12777,s12778,s12779,s12780,s12781,s12782,s12783,s12784,s12785,s12786,s12787,s12788,s12789,s12790,s12791,s12792,s12793,s12794,s12795,s12796,s12797,s12798,s12799,

s12800,s12801,s12802,s12803,s12804,s12805,s12806,s12807,s12808,s12809,s12810,s12811,s12812,s12813,s12814,s12815,s12816,s12817,s12818,s12819,s12820,s12821,s12822,s12823,s12824,s12825,s12826,s12827,s12828,s12829,s12830,s12831,s12832,s12833,s12834,s12835,s12836,s12837,s12838,s12839,s12840,s12841,s12842,s12843,s12844,s12845,s12846,s12847,s12848,s12849,s12850,s12851,s12852,s12853,s12854,s12855,s12856,s12857,s12858,s12859,s12860,s12861,s12862,s12863,s12864,s12865,s12866,s12867,s12868,s12869,s12870,s12871,s12872,s12873,s12874,s12875,s12876,s12877,s12878,s12879,

s12880,s12881,s12882,s12883,s12884,s12885,s12886,s12887,s12888,s12889,s12890,s12891,s12892,s12893,s12894,s12895,s12896,s12897,s12898,s12899,s12900,s12901,s12902,s12903,s12904,s12905,s12906,s12907,s12908,s12909,s12910,s12911,s12912,s12913,s12914,s12915,s12916,s12917,s12918,s12919,s12920,s12921,s12922,s12923,s12924,s12925,s12926,s12927,s12928,s12929,s12930,s12931,s12932,s12933,s12934,s12935,s12936,s12937,s12938,s12939,s12940,s12941,s12942,s12943,s12944,s12945,s12946,s12947,s12948,s12949,s12950,s12951,s12952,s12953,s12954,s12955,s12956,s12957,s12958,s12959,

s12960,s12961,s12962,s12963,s12964,s12965,s12966,s12967,s12968,s12969,s12970,s12971,s12972,s12973,s12974,s12975,s12976,s12977,s12978,s12979,s12980,s12981,s12982,s12983,s12984,s12985,s12986,s12987,s12988,s12989,s12990,s12991,s12992,s12993,s12994,s12995,s12996,s12997,s12998,s12999,s13000,s13001,s13002,s13003,s13004,s13005,s13006,s13007,s13008,s13009,s13010,s13011,s13012,s13013,s13014,s13015,s13016,s13017,s13018,s13019,s13020,s13021,s13022,s13023,s13024,s13025,s13026,s13027,s13028,s13029,s13030,s13031,s13032,s13033,s13034,s13035,s13036,s13037,s13038,s13039,

s13040,s13041,s13042,s13043,s13044,s13045,s13046,s13047,s13048,s13049,s13050,s13051,s13052,s13053,s13054,s13055,s13056,s13057,s13058,s13059,s13060,s13061,s13062,s13063,s13064,s13065,s13066,s13067,s13068,s13069,s13070,s13071,s13072,s13073,s13074,s13075,s13076,s13077,s13078,s13079,s13080,s13081,s13082,s13083,s13084,s13085,s13086,s13087,s13088,s13089,s13090,s13091,s13092,s13093,s13094,s13095,s13096,s13097,s13098,s13099,s13100,s13101,s13102,s13103,s13104,s13105,s13106,s13107,s13108,s13109,s13110,s13111,s13112,s13113,s13114,s13115,s13116,s13117,s13118,s13119,

s13120,s13121,s13122,s13123,s13124,s13125,s13126,s13127,s13128,s13129,s13130,s13131,s13132,s13133,s13134,s13135,s13136,s13137,s13138,s13139,s13140,s13141,s13142,s13143,s13144,s13145,s13146,s13147,s13148,s13149,s13150,s13151,s13152,s13153,s13154,s13155,s13156,s13157,s13158,s13159,s13160,s13161,s13162,s13163,s13164,s13165,s13166,s13167,s13168,s13169,s13170,s13171,s13172,s13173,s13174,s13175,s13176,s13177,s13178,s13179,s13180,s13181,s13182,s13183,s13184,s13185,s13186,s13187,s13188,s13189,s13190,s13191,s13192,s13193,s13194,s13195,s13196,s13197,s13198,s13199,

s13200,s13201,s13202,s13203,s13204,s13205,s13206,s13207,s13208,s13209,s13210,s13211,s13212,s13213,s13214,s13215,s13216,s13217,s13218,s13219,s13220,s13221,s13222,s13223,s13224,s13225,s13226,s13227,s13228,s13229,s13230,s13231,s13232,s13233,s13234,s13235,s13236,s13237,s13238,s13239,s13240,s13241,s13242,s13243,s13244,s13245,s13246,s13247,s13248,s13249,s13250,s13251,s13252,s13253,s13254,s13255,s13256,s13257,s13258,s13259,s13260,s13261,s13262,s13263,s13264,s13265,s13266,s13267,s13268,s13269,s13270,s13271,s13272,s13273,s13274,s13275,s13276,s13277,s13278,s13279,

s13280,s13281,s13282,s13283,s13284,s13285,s13286,s13287,s13288,s13289,s13290,s13291,s13292,s13293,s13294,s13295,s13296,s13297,s13298,s13299,s13300,s13301,s13302,s13303,s13304,s13305,s13306,s13307,s13308,s13309,s13310,s13311,s13312,s13313,s13314,s13315,s13316,s13317,s13318,s13319,s13320,s13321,s13322,s13323,s13324,s13325,s13326,s13327,s13328,s13329,s13330,s13331,s13332,s13333,s13334,s13335,s13336,s13337,s13338,s13339,s13340,s13341,s13342,s13343,s13344,s13345,s13346,s13347,s13348,s13349,s13350,s13351,s13352,s13353,s13354,s13355,s13356,s13357,s13358,s13359,

s13360,s13361,s13362,s13363,s13364,s13365,s13366,s13367,s13368,s13369,s13370,s13371,s13372,s13373,s13374,s13375,s13376,s13377,s13378,s13379,s13380,s13381,s13382,s13383,s13384,s13385,s13386,s13387,s13388,s13389,s13390,s13391,s13392,s13393,s13394,s13395,s13396,s13397,s13398,s13399,s13400,s13401,s13402,s13403,s13404,s13405,s13406,s13407,s13408,s13409,s13410,s13411,s13412,s13413,s13414,s13415,s13416,s13417,s13418,s13419,s13420,s13421,s13422,s13423,s13424,s13425,s13426,s13427,s13428,s13429,s13430,s13431,s13432,s13433,s13434,s13435,s13436,s13437,s13438,s13439,

s13440,s13441,s13442,s13443,s13444,s13445,s13446,s13447,s13448,s13449,s13450,s13451,s13452,s13453,s13454,s13455,s13456,s13457,s13458,s13459,s13460,s13461,s13462,s13463,s13464,s13465,s13466,s13467,s13468,s13469,s13470,s13471,s13472,s13473,s13474,s13475,s13476,s13477,s13478,s13479,s13480,s13481,s13482,s13483,s13484,s13485,s13486,s13487,s13488,s13489,s13490,s13491,s13492,s13493,s13494,s13495,s13496,s13497,s13498,s13499,s13500,s13501,s13502,s13503,s13504,s13505,s13506,s13507,s13508,s13509,s13510,s13511,s13512,s13513,s13514,s13515,s13516,s13517,s13518,s13519,

s13520,s13521,s13522,s13523,s13524,s13525,s13526,s13527,s13528,s13529,s13530,s13531,s13532,s13533,s13534,s13535,s13536,s13537,s13538,s13539,s13540,s13541,s13542,s13543,s13544,s13545,s13546,s13547,s13548,s13549,s13550,s13551,s13552,s13553,s13554,s13555,s13556,s13557,s13558,s13559,s13560,s13561,s13562,s13563,s13564,s13565,s13566,s13567,s13568,s13569,s13570,s13571,s13572,s13573,s13574,s13575,s13576,s13577,s13578,s13579,s13580,s13581,s13582,s13583,s13584,s13585,s13586,s13587,s13588,s13589,s13590,s13591,s13592,s13593,s13594,s13595,s13596,s13597,s13598,s13599,

s13600,s13601,s13602,s13603,s13604,s13605,s13606,s13607,s13608,s13609,s13610,s13611,s13612,s13613,s13614,s13615,s13616,s13617,s13618,s13619,s13620,s13621,s13622,s13623,s13624,s13625,s13626,s13627,s13628,s13629,s13630,s13631,s13632,s13633,s13634,s13635,s13636,s13637,s13638,s13639,s13640,s13641,s13642,s13643,s13644,s13645,s13646,s13647,s13648,s13649,s13650,s13651,s13652,s13653,s13654,s13655,s13656,s13657,s13658,s13659,s13660,s13661,s13662,s13663,s13664,s13665,s13666,s13667,s13668,s13669,s13670,s13671,s13672,s13673,s13674,s13675,s13676,s13677,s13678,s13679,

s13680,s13681,s13682,s13683,s13684,s13685,s13686,s13687,s13688,s13689,s13690,s13691,s13692,s13693,s13694,s13695,s13696,s13697,s13698,s13699,s13700,s13701,s13702,s13703,s13704,s13705,s13706,s13707,s13708,s13709,s13710,s13711,s13712,s13713,s13714,s13715,s13716,s13717,s13718,s13719,s13720,s13721,s13722,s13723,s13724,s13725,s13726,s13727,s13728,s13729,s13730,s13731,s13732,s13733,s13734,s13735,s13736,s13737,s13738,s13739,s13740,s13741,s13742,s13743,s13744,s13745,s13746,s13747,s13748,s13749,s13750,s13751,s13752,s13753,s13754,s13755,s13756,s13757,s13758,s13759,

s13760,s13761,s13762,s13763,s13764,s13765,s13766,s13767,s13768,s13769,s13770,s13771,s13772,s13773,s13774,s13775,s13776,s13777,s13778,s13779,s13780,s13781,s13782,s13783,s13784,s13785,s13786,s13787,s13788,s13789,s13790,s13791,s13792,s13793,s13794,s13795,s13796,s13797,s13798,s13799,s13800,s13801,s13802,s13803,s13804,s13805,s13806,s13807,s13808,s13809,s13810,s13811,s13812,s13813,s13814,s13815,s13816,s13817,s13818,s13819,s13820,s13821,s13822,s13823,s13824,s13825,s13826,s13827,s13828,s13829,s13830,s13831,s13832,s13833,s13834,s13835,s13836,s13837,s13838,s13839,

s13840,s13841,s13842,s13843,s13844,s13845,s13846,s13847,s13848,s13849,s13850,s13851,s13852,s13853,s13854,s13855,s13856,s13857,s13858,s13859,s13860,s13861,s13862,s13863,s13864,s13865,s13866,s13867,s13868,s13869,s13870,s13871,s13872,s13873,s13874,s13875,s13876,s13877,s13878,s13879,s13880,s13881,s13882,s13883,s13884,s13885,s13886,s13887,s13888,s13889,s13890,s13891,s13892,s13893,s13894,s13895,s13896,s13897,s13898,s13899,s13900,s13901,s13902,s13903,s13904,s13905,s13906,s13907,s13908,s13909,s13910,s13911,s13912,s13913,s13914,s13915,s13916,s13917,s13918,s13919,

s13920,s13921,s13922,s13923,s13924,s13925,s13926,s13927,s13928,s13929,s13930,s13931,s13932,s13933,s13934,s13935,s13936,s13937,s13938,s13939,s13940,s13941,s13942,s13943,s13944,s13945,s13946,s13947,s13948,s13949,s13950,s13951,s13952,s13953,s13954,s13955,s13956,s13957,s13958,s13959,s13960,s13961,s13962,s13963,s13964,s13965,s13966,s13967,s13968,s13969,s13970,s13971,s13972,s13973,s13974,s13975,s13976,s13977,s13978,s13979,s13980,s13981,s13982,s13983,s13984,s13985,s13986,s13987,s13988,s13989,s13990,s13991,s13992,s13993,s13994,s13995,s13996,s13997,s13998,s13999,

s14000,s14001,s14002,s14003,s14004,s14005,s14006,s14007,s14008,s14009,s14010,s14011,s14012,s14013,s14014,s14015,s14016,s14017,s14018,s14019,s14020,s14021,s14022,s14023,s14024,s14025,s14026,s14027,s14028,s14029,s14030,s14031,s14032,s14033,s14034,s14035,s14036,s14037,s14038,s14039,s14040,s14041,s14042,s14043,s14044,s14045,s14046,s14047,s14048,s14049,s14050,s14051,s14052,s14053,s14054,s14055,s14056,s14057,s14058,s14059,s14060,s14061,s14062,s14063,s14064,s14065,s14066,s14067,s14068,s14069,s14070,s14071,s14072,s14073,s14074,s14075,s14076,s14077,s14078,s14079,

s14080,s14081,s14082,s14083,s14084,s14085,s14086,s14087,s14088,s14089,s14090,s14091,s14092,s14093,s14094,s14095,s14096,s14097,s14098,s14099,s14100,s14101,s14102,s14103,s14104,s14105,s14106,s14107,s14108,s14109,s14110,s14111,s14112,s14113,s14114,s14115,s14116,s14117,s14118,s14119,s14120,s14121,s14122,s14123,s14124,s14125,s14126,s14127,s14128,s14129,s14130,s14131,s14132,s14133,s14134,s14135,s14136,s14137,s14138,s14139,s14140,s14141,s14142,s14143,s14144,s14145,s14146,s14147,s14148,s14149,s14150,s14151,s14152,s14153,s14154,s14155,s14156,s14157,s14158,s14159,

s14160,s14161,s14162,s14163,s14164,s14165,s14166,s14167,s14168,s14169,s14170,s14171,s14172,s14173,s14174,s14175,s14176,s14177,s14178,s14179,s14180,s14181,s14182,s14183,s14184,s14185,s14186,s14187,s14188,s14189,s14190,s14191,s14192,s14193,s14194,s14195,s14196,s14197,s14198,s14199,s14200,s14201,s14202,s14203,s14204,s14205,s14206,s14207,s14208,s14209,s14210,s14211,s14212,s14213,s14214,s14215,s14216,s14217,s14218,s14219,s14220,s14221,s14222,s14223,s14224,s14225,s14226,s14227,s14228,s14229,s14230,s14231,s14232,s14233,s14234,s14235,s14236,s14237,s14238,s14239,

s14240,s14241,s14242,s14243,s14244,s14245,s14246,s14247,s14248,s14249,s14250,s14251,s14252,s14253,s14254,s14255,s14256,s14257,s14258,s14259,s14260,s14261,s14262,s14263,s14264,s14265,s14266,s14267,s14268,s14269,s14270,s14271,s14272,s14273,s14274,s14275,s14276,s14277,s14278,s14279,s14280,s14281,s14282,s14283,s14284,s14285,s14286,s14287,s14288,s14289,s14290,s14291,s14292,s14293,s14294,s14295,s14296,s14297,s14298,s14299,s14300,s14301,s14302,s14303,s14304,s14305,s14306,s14307,s14308,s14309,s14310,s14311,s14312,s14313,s14314,s14315,s14316,s14317,s14318,s14319,

s14320,s14321,s14322,s14323,s14324,s14325,s14326,s14327,s14328,s14329,s14330,s14331,s14332,s14333,s14334,s14335,s14336,s14337,s14338,s14339,s14340,s14341,s14342,s14343,s14344,s14345,s14346,s14347,s14348,s14349,s14350,s14351,s14352,s14353,s14354,s14355,s14356,s14357,s14358,s14359,s14360,s14361,s14362,s14363,s14364,s14365,s14366,s14367,s14368,s14369,s14370,s14371,s14372,s14373,s14374,s14375,s14376,s14377,s14378,s14379,s14380,s14381,s14382,s14383,s14384,s14385,s14386,s14387,s14388,s14389,s14390,s14391,s14392,s14393,s14394,s14395,s14396,s14397,s14398,s14399,

s14400,s14401,s14402,s14403,s14404,s14405,s14406,s14407,s14408,s14409,s14410,s14411,s14412,s14413,s14414,s14415,s14416,s14417,s14418,s14419,s14420,s14421,s14422,s14423,s14424,s14425,s14426,s14427,s14428,s14429,s14430,s14431,s14432,s14433,s14434,s14435,s14436,s14437,s14438,s14439,s14440,s14441,s14442,s14443,s14444,s14445,s14446,s14447,s14448,s14449,s14450,s14451,s14452,s14453,s14454,s14455,s14456,s14457,s14458,s14459,s14460,s14461,s14462,s14463,s14464,s14465,s14466,s14467,s14468,s14469,s14470,s14471,s14472,s14473,s14474,s14475,s14476,s14477,s14478,s14479,

s14480,s14481,s14482,s14483,s14484,s14485,s14486,s14487,s14488,s14489,s14490,s14491,s14492,s14493,s14494,s14495,s14496,s14497,s14498,s14499,s14500,s14501,s14502,s14503,s14504,s14505,s14506,s14507,s14508,s14509,s14510,s14511,s14512,s14513,s14514,s14515,s14516,s14517,s14518,s14519,s14520,s14521,s14522,s14523,s14524,s14525,s14526,s14527,s14528,s14529,s14530,s14531,s14532,s14533,s14534,s14535,s14536,s14537,s14538,s14539,s14540,s14541,s14542,s14543,s14544,s14545,s14546,s14547,s14548,s14549,s14550,s14551,s14552,s14553,s14554,s14555,s14556,s14557,s14558,s14559,

s14560,s14561,s14562,s14563,s14564,s14565,s14566,s14567,s14568,s14569,s14570,s14571,s14572,s14573,s14574,s14575,s14576,s14577,s14578,s14579,s14580,s14581,s14582,s14583,s14584,s14585,s14586,s14587,s14588,s14589,s14590,s14591,s14592,s14593,s14594,s14595,s14596,s14597,s14598,s14599,s14600,s14601,s14602,s14603,s14604,s14605,s14606,s14607,s14608,s14609,s14610,s14611,s14612,s14613,s14614,s14615,s14616,s14617,s14618,s14619,s14620,s14621,s14622,s14623,s14624,s14625,s14626,s14627,s14628,s14629,s14630,s14631,s14632,s14633,s14634,s14635,s14636,s14637,s14638,s14639,

s14640,s14641,s14642,s14643,s14644,s14645,s14646,s14647,s14648,s14649,s14650,s14651,s14652,s14653,s14654,s14655,s14656,s14657,s14658,s14659,s14660,s14661,s14662,s14663,s14664,s14665,s14666,s14667,s14668,s14669,s14670,s14671,s14672,s14673,s14674,s14675,s14676,s14677,s14678,s14679,s14680,s14681,s14682,s14683,s14684,s14685,s14686,s14687,s14688,s14689,s14690,s14691,s14692,s14693,s14694,s14695,s14696,s14697,s14698,s14699,s14700,s14701,s14702,s14703,s14704,s14705,s14706,s14707,s14708,s14709,s14710,s14711,s14712,s14713,s14714,s14715,s14716,s14717,s14718,s14719,

s14720,s14721,s14722,s14723,s14724,s14725,s14726,s14727,s14728,s14729,s14730,s14731,s14732,s14733,s14734,s14735,s14736,s14737,s14738,s14739,s14740,s14741,s14742,s14743,s14744,s14745,s14746,s14747,s14748,s14749,s14750,s14751,s14752,s14753,s14754,s14755,s14756,s14757,s14758,s14759,s14760,s14761,s14762,s14763,s14764,s14765,s14766,s14767,s14768,s14769,s14770,s14771,s14772,s14773,s14774,s14775,s14776,s14777,s14778,s14779,s14780,s14781,s14782,s14783,s14784,s14785,s14786,s14787,s14788,s14789,s14790,s14791,s14792,s14793,s14794,s14795,s14796,s14797,s14798,s14799,

s14800,s14801,s14802,s14803,s14804,s14805,s14806,s14807,s14808,s14809,s14810,s14811,s14812,s14813,s14814,s14815,s14816,s14817,s14818,s14819,s14820,s14821,s14822,s14823,s14824,s14825,s14826,s14827,s14828,s14829,s14830,s14831,s14832,s14833,s14834,s14835,s14836,s14837,s14838,s14839,s14840,s14841,s14842,s14843,s14844,s14845,s14846,s14847,s14848,s14849,s14850,s14851,s14852,s14853,s14854,s14855,s14856,s14857,s14858,s14859,s14860,s14861,s14862,s14863,s14864,s14865,s14866,s14867,s14868,s14869,s14870,s14871,s14872,s14873,s14874,s14875,s14876,s14877,s14878,s14879,

s14880,s14881,s14882,s14883,s14884,s14885,s14886,s14887,s14888,s14889,s14890,s14891,s14892,s14893,s14894,s14895,s14896,s14897,s14898,s14899,s14900,s14901,s14902,s14903,s14904,s14905,s14906,s14907,s14908,s14909,s14910,s14911,s14912,s14913,s14914,s14915,s14916,s14917,s14918,s14919,s14920,s14921,s14922,s14923,s14924,s14925,s14926,s14927,s14928,s14929,s14930,s14931,s14932,s14933,s14934,s14935,s14936,s14937,s14938,s14939,s14940,s14941,s14942,s14943,s14944,s14945,s14946,s14947,s14948,s14949,s14950,s14951,s14952,s14953,s14954,s14955,s14956,s14957,s14958,s14959,

s14960,s14961,s14962,s14963,s14964,s14965,s14966,s14967,s14968,s14969,s14970,s14971,s14972,s14973,s14974,s14975,s14976,s14977,s14978,s14979,s14980,s14981,s14982,s14983,s14984,s14985,s14986,s14987,s14988,s14989,s14990,s14991,s14992,s14993,s14994,s14995,s14996,s14997,s14998,s14999,s15000,s15001,s15002,s15003,s15004,s15005,s15006,s15007,s15008,s15009,s15010,s15011,s15012,s15013,s15014,s15015,s15016,s15017,s15018,s15019,s15020,s15021,s15022,s15023,s15024,s15025,s15026,s15027,s15028,s15029,s15030,s15031,s15032,s15033,s15034,s15035,s15036,s15037,s15038,s15039,

s15040,s15041,s15042,s15043,s15044,s15045,s15046,s15047,s15048,s15049,s15050,s15051,s15052,s15053,s15054,s15055,s15056,s15057,s15058,s15059,s15060,s15061,s15062,s15063,s15064,s15065,s15066,s15067,s15068,s15069,s15070,s15071,s15072,s15073,s15074,s15075,s15076,s15077,s15078,s15079,s15080,s15081,s15082,s15083,s15084,s15085,s15086,s15087,s15088,s15089,s15090,s15091,s15092,s15093,s15094,s15095,s15096,s15097,s15098,s15099,s15100,s15101,s15102,s15103,s15104,s15105,s15106,s15107,s15108,s15109,s15110,s15111,s15112,s15113,s15114,s15115,s15116,s15117,s15118,s15119,

s15120,s15121,s15122,s15123,s15124,s15125,s15126,s15127,s15128,s15129,s15130,s15131,s15132,s15133,s15134,s15135,s15136,s15137,s15138,s15139,s15140,s15141,s15142,s15143,s15144,s15145,s15146,s15147,s15148,s15149,s15150,s15151,s15152,s15153,s15154,s15155,s15156,s15157,s15158,s15159,s15160,s15161,s15162,s15163,s15164,s15165,s15166,s15167,s15168,s15169,s15170,s15171,s15172,s15173,s15174,s15175,s15176,s15177,s15178,s15179,s15180,s15181,s15182,s15183,s15184,s15185,s15186,s15187,s15188,s15189,s15190,s15191,s15192,s15193,s15194,s15195,s15196,s15197,s15198,s15199,

s15200,s15201,s15202,s15203,s15204,s15205,s15206,s15207,s15208,s15209,s15210,s15211,s15212,s15213,s15214,s15215,s15216,s15217,s15218,s15219,s15220,s15221,s15222,s15223,s15224,s15225,s15226,s15227,s15228,s15229,s15230,s15231,s15232,s15233,s15234,s15235,s15236,s15237,s15238,s15239,s15240,s15241,s15242,s15243,s15244,s15245,s15246,s15247,s15248,s15249,s15250,s15251,s15252,s15253,s15254,s15255,s15256,s15257,s15258,s15259,s15260,s15261,s15262,s15263,s15264,s15265,s15266,s15267,s15268,s15269,s15270,s15271,s15272,s15273,s15274,s15275,s15276,s15277,s15278,s15279,

s15280,s15281,s15282,s15283,s15284,s15285,s15286,s15287,s15288,s15289,s15290,s15291,s15292,s15293,s15294,s15295,s15296,s15297,s15298,s15299,s15300,s15301,s15302,s15303,s15304,s15305,s15306,s15307,s15308,s15309,s15310,s15311,s15312,s15313,s15314,s15315,s15316,s15317,s15318,s15319,s15320,s15321,s15322,s15323,s15324,s15325,s15326,s15327,s15328,s15329,s15330,s15331,s15332,s15333,s15334,s15335,s15336,s15337,s15338,s15339,s15340,s15341,s15342,s15343,s15344,s15345,s15346,s15347,s15348,s15349,s15350,s15351,s15352,s15353,s15354,s15355,s15356,s15357,s15358,s15359,

s15360,s15361,s15362,s15363,s15364,s15365,s15366,s15367,s15368,s15369,s15370,s15371,s15372,s15373,s15374,s15375,s15376,s15377,s15378,s15379,s15380,s15381,s15382,s15383,s15384,s15385,s15386,s15387,s15388,s15389,s15390,s15391,s15392,s15393,s15394,s15395,s15396,s15397,s15398,s15399,s15400,s15401,s15402,s15403,s15404,s15405,s15406,s15407,s15408,s15409,s15410,s15411,s15412,s15413,s15414,s15415,s15416,s15417,s15418,s15419,s15420,s15421,s15422,s15423,s15424,s15425,s15426,s15427,s15428,s15429,s15430,s15431,s15432,s15433,s15434,s15435,s15436,s15437,s15438,s15439,

s15440,s15441,s15442,s15443,s15444,s15445,s15446,s15447,s15448,s15449,s15450,s15451,s15452,s15453,s15454,s15455,s15456,s15457,s15458,s15459,s15460,s15461,s15462,s15463,s15464,s15465,s15466,s15467,s15468,s15469,s15470,s15471,s15472,s15473,s15474,s15475,s15476,s15477,s15478,s15479,s15480,s15481,s15482,s15483,s15484,s15485,s15486,s15487,s15488,s15489,s15490,s15491,s15492,s15493,s15494,s15495,s15496,s15497,s15498,s15499,s15500,s15501,s15502,s15503,s15504,s15505,s15506,s15507,s15508,s15509,s15510,s15511,s15512,s15513,s15514,s15515,s15516,s15517,s15518,s15519,

s15520,s15521,s15522,s15523,s15524,s15525,s15526,s15527,s15528,s15529,s15530,s15531,s15532,s15533,s15534,s15535,s15536,s15537,s15538,s15539,s15540,s15541,s15542,s15543,s15544,s15545,s15546,s15547,s15548,s15549,s15550,s15551,s15552,s15553,s15554,s15555,s15556,s15557,s15558,s15559,s15560,s15561,s15562,s15563,s15564,s15565,s15566,s15567,s15568,s15569,s15570,s15571,s15572,s15573,s15574,s15575,s15576,s15577,s15578,s15579,s15580,s15581,s15582,s15583,s15584,s15585,s15586,s15587,s15588,s15589,s15590,s15591,s15592,s15593,s15594,s15595,s15596,s15597,s15598,s15599,

s15600,s15601,s15602,s15603,s15604,s15605,s15606,s15607,s15608,s15609,s15610,s15611,s15612,s15613,s15614,s15615,s15616,s15617,s15618,s15619,s15620,s15621,s15622,s15623,s15624,s15625,s15626,s15627,s15628,s15629,s15630,s15631,s15632,s15633,s15634,s15635,s15636,s15637,s15638,s15639,s15640,s15641,s15642,s15643,s15644,s15645,s15646,s15647,s15648,s15649,s15650,s15651,s15652,s15653,s15654,s15655,s15656,s15657,s15658,s15659,s15660,s15661,s15662,s15663,s15664,s15665,s15666,s15667,s15668,s15669,s15670,s15671,s15672,s15673,s15674,s15675,s15676,s15677,s15678,s15679,

s15680,s15681,s15682,s15683,s15684,s15685,s15686,s15687,s15688,s15689,s15690,s15691,s15692,s15693,s15694,s15695,s15696,s15697,s15698,s15699,s15700,s15701,s15702,s15703,s15704,s15705,s15706,s15707,s15708,s15709,s15710,s15711,s15712,s15713,s15714,s15715,s15716,s15717,s15718,s15719,s15720,s15721,s15722,s15723,s15724,s15725,s15726,s15727,s15728,s15729,s15730,s15731,s15732,s15733,s15734,s15735,s15736,s15737,s15738,s15739,s15740,s15741,s15742,s15743,s15744,s15745,s15746,s15747,s15748,s15749,s15750,s15751,s15752,s15753,s15754,s15755,s15756,s15757,s15758,s15759,

s15760,s15761,s15762,s15763,s15764,s15765,s15766,s15767,s15768,s15769,s15770,s15771,s15772,s15773,s15774,s15775,s15776,s15777,s15778,s15779,s15780,s15781,s15782,s15783,s15784,s15785,s15786,s15787,s15788,s15789,s15790,s15791,s15792,s15793,s15794,s15795,s15796,s15797,s15798,s15799,s15800,s15801,s15802,s15803,s15804,s15805,s15806,s15807,s15808,s15809,s15810,s15811,s15812,s15813,s15814,s15815,s15816,s15817,s15818,s15819,s15820,s15821,s15822,s15823,s15824,s15825,s15826,s15827,s15828,s15829,s15830,s15831,s15832,s15833,s15834,s15835,s15836,s15837,s15838,s15839,

s15840,s15841,s15842,s15843,s15844,s15845,s15846,s15847,s15848,s15849,s15850,s15851,s15852,s15853,s15854,s15855,s15856,s15857,s15858,s15859,s15860,s15861,s15862,s15863,s15864,s15865,s15866,s15867,s15868,s15869,s15870,s15871,s15872,s15873,s15874,s15875,s15876,s15877,s15878,s15879,s15880,s15881,s15882,s15883,s15884,s15885,s15886,s15887,s15888,s15889,s15890,s15891,s15892,s15893,s15894,s15895,s15896,s15897,s15898,s15899,s15900,s15901,s15902,s15903,s15904,s15905,s15906,s15907,s15908,s15909,s15910,s15911,s15912,s15913,s15914,s15915,s15916,s15917,s15918,s15919,

s15920,s15921,s15922,s15923,s15924,s15925,s15926,s15927,s15928,s15929,s15930,s15931,s15932,s15933,s15934,s15935,s15936,s15937,s15938,s15939,s15940,s15941,s15942,s15943,s15944,s15945,s15946,s15947,s15948,s15949,s15950,s15951,s15952,s15953,s15954,s15955,s15956,s15957,s15958,s15959,s15960,s15961,s15962,s15963,s15964,s15965,s15966,s15967,s15968,s15969,s15970,s15971,s15972,s15973,s15974,s15975,s15976,s15977,s15978,s15979,s15980,s15981,s15982,s15983,s15984,s15985,s15986,s15987,s15988,s15989,s15990,s15991,s15992,s15993,s15994,s15995,s15996,s15997,s15998,s15999,

s16000,s16001,s16002,s16003,s16004,s16005,s16006,s16007,s16008,s16009,s16010,s16011,s16012,s16013,s16014,s16015,s16016,s16017,s16018,s16019,s16020,s16021,s16022,s16023,s16024,s16025,s16026,s16027,s16028,s16029,s16030,s16031,s16032,s16033,s16034,s16035,s16036,s16037,s16038,s16039,s16040,s16041,s16042,s16043,s16044,s16045,s16046,s16047,s16048,s16049,s16050,s16051,s16052,s16053,s16054,s16055,s16056,s16057,s16058,s16059,s16060,s16061,s16062,s16063,s16064,s16065,s16066,s16067,s16068,s16069,s16070,s16071,s16072,s16073,s16074,s16075,s16076,s16077,s16078,s16079,

s16080,s16081,s16082,s16083,s16084,s16085,s16086,s16087,s16088,s16089,s16090,s16091,s16092,s16093,s16094,s16095,s16096,s16097,s16098,s16099,s16100,s16101,s16102,s16103,s16104,s16105,s16106,s16107,s16108,s16109,s16110,s16111,s16112,s16113,s16114,s16115,s16116,s16117,s16118,s16119,s16120,s16121,s16122,s16123,s16124,s16125,s16126,s16127,s16128,s16129,s16130,s16131,s16132,s16133,s16134,s16135,s16136,s16137,s16138,s16139,s16140,s16141,s16142,s16143,s16144,s16145,s16146,s16147,s16148,s16149,s16150,s16151,s16152,s16153,s16154,s16155,s16156,s16157,s16158,s16159,

s16160,s16161,s16162,s16163,s16164,s16165,s16166,s16167,s16168,s16169,s16170,s16171,s16172,s16173,s16174,s16175,s16176,s16177,s16178,s16179,s16180,s16181,s16182,s16183,s16184,s16185,s16186,s16187,s16188,s16189,s16190,s16191,s16192,s16193,s16194,s16195,s16196,s16197,s16198,s16199,s16200,s16201,s16202,s16203,s16204,s16205,s16206,s16207,s16208,s16209,s16210,s16211,s16212,s16213,s16214,s16215,s16216,s16217,s16218,s16219,s16220,s16221,s16222,s16223,s16224,s16225,s16226,s16227,s16228,s16229,s16230,s16231,s16232,s16233,s16234,s16235,s16236,s16237,s16238,s16239,

s16240,s16241,s16242,s16243,s16244,s16245,s16246,s16247,s16248,s16249,s16250,s16251,s16252,s16253,s16254,s16255,s16256,s16257,s16258,s16259,s16260,s16261,s16262,s16263,s16264,s16265,s16266,s16267,s16268,s16269,s16270,s16271,s16272,s16273,s16274,s16275,s16276,s16277,s16278,s16279,s16280,s16281,s16282,s16283,s16284,s16285,s16286,s16287,s16288,s16289,s16290,s16291,s16292,s16293,s16294,s16295,s16296,s16297,s16298,s16299,s16300,s16301,s16302,s16303,s16304,s16305,s16306,s16307,s16308,s16309,s16310,s16311,s16312,s16313,s16314,s16315,s16316,s16317,s16318,s16319,

s16320,s16321,s16322,s16323,s16324,s16325,s16326,s16327,s16328,s16329,s16330,s16331,s16332,s16333,s16334,s16335,s16336,s16337,s16338,s16339,s16340,s16341,s16342,s16343,s16344,s16345,s16346,s16347,s16348,s16349,s16350,s16351,s16352,s16353,s16354,s16355,s16356,s16357,s16358,s16359,s16360,s16361,s16362,s16363,s16364,s16365,s16366,s16367,s16368,s16369,s16370,s16371,s16372,s16373,s16374,s16375,s16376,s16377,s16378,s16379,s16380,s16381,s16382,s16383,s16384,s16385,s16386,s16387,s16388,s16389,s16390,s16391,s16392,s16393,s16394,s16395,s16396,s16397,s16398,s16399,

s16400,s16401,s16402,s16403,s16404,s16405,s16406,s16407,s16408,s16409,s16410,s16411,s16412,s16413,s16414,s16415,s16416,s16417,s16418,s16419,s16420,s16421,s16422,s16423,s16424,s16425,s16426,s16427,s16428,s16429,s16430,s16431,s16432,s16433,s16434,s16435,s16436,s16437,s16438,s16439,s16440,s16441,s16442,s16443,s16444,s16445,s16446,s16447,s16448,s16449,s16450,s16451,s16452,s16453,s16454,s16455,s16456,s16457,s16458,s16459,s16460,s16461,s16462,s16463,s16464,s16465,s16466,s16467,s16468,s16469,s16470,s16471,s16472,s16473,s16474,s16475,s16476,s16477,s16478,s16479,

s16480,s16481,s16482,s16483,s16484,s16485,s16486,s16487,s16488,s16489,s16490,s16491,s16492,s16493,s16494,s16495,s16496,s16497,s16498,s16499,s16500,s16501,s16502,s16503,s16504,s16505,s16506,s16507,s16508,s16509,s16510,s16511,s16512,s16513,s16514,s16515,s16516,s16517,s16518,s16519,s16520,s16521,s16522,s16523,s16524,s16525,s16526,s16527,s16528,s16529,s16530,s16531,s16532,s16533,s16534,s16535,s16536,s16537,s16538,s16539,s16540,s16541,s16542,s16543,s16544,s16545,s16546,s16547,s16548,s16549,s16550,s16551,s16552,s16553,s16554,s16555,s16556,s16557,s16558,s16559,

s16560,s16561,s16562,s16563,s16564,s16565,s16566,s16567,s16568,s16569,s16570,s16571,s16572,s16573,s16574,s16575,s16576,s16577,s16578,s16579,s16580,s16581,s16582,s16583,s16584,s16585,s16586,s16587,s16588,s16589,s16590,s16591,s16592,s16593,s16594,s16595,s16596,s16597,s16598,s16599,s16600,s16601,s16602,s16603,s16604,s16605,s16606,s16607,s16608,s16609,s16610,s16611,s16612,s16613,s16614,s16615,s16616,s16617,s16618,s16619,s16620,s16621,s16622,s16623,s16624,s16625,s16626,s16627,s16628,s16629,s16630,s16631,s16632,s16633,s16634,s16635,s16636,s16637,s16638,s16639,

s16640,s16641,s16642,s16643,s16644,s16645,s16646,s16647,s16648,s16649,s16650,s16651,s16652,s16653,s16654,s16655,s16656,s16657,s16658,s16659,s16660,s16661,s16662,s16663,s16664,s16665,s16666,s16667,s16668,s16669,s16670,s16671,s16672,s16673,s16674,s16675,s16676,s16677,s16678,s16679,s16680,s16681,s16682,s16683,s16684,s16685,s16686,s16687,s16688,s16689,s16690,s16691,s16692,s16693,s16694,s16695,s16696,s16697,s16698,s16699,s16700,s16701,s16702,s16703,s16704,s16705,s16706,s16707,s16708,s16709,s16710,s16711,s16712,s16713,s16714,s16715,s16716,s16717,s16718,s16719,

s16720,s16721,s16722,s16723,s16724,s16725,s16726,s16727,s16728,s16729,s16730,s16731,s16732,s16733,s16734,s16735,s16736,s16737,s16738,s16739,s16740,s16741,s16742,s16743,s16744,s16745,s16746,s16747,s16748,s16749,s16750,s16751,s16752,s16753,s16754,s16755,s16756,s16757,s16758,s16759,s16760,s16761,s16762,s16763,s16764,s16765,s16766,s16767,s16768,s16769,s16770,s16771,s16772,s16773,s16774,s16775,s16776,s16777,s16778,s16779,s16780,s16781,s16782,s16783,s16784,s16785,s16786,s16787,s16788,s16789,s16790,s16791,s16792,s16793,s16794,s16795,s16796,s16797,s16798,s16799,

s16800,s16801,s16802,s16803,s16804,s16805,s16806,s16807,s16808,s16809,s16810,s16811,s16812,s16813,s16814,s16815,s16816,s16817,s16818,s16819,s16820,s16821,s16822,s16823,s16824,s16825,s16826,s16827,s16828,s16829,s16830,s16831,s16832,s16833,s16834,s16835,s16836,s16837,s16838,s16839,s16840,s16841,s16842,s16843,s16844,s16845,s16846,s16847,s16848,s16849,s16850,s16851,s16852,s16853,s16854,s16855,s16856,s16857,s16858,s16859,s16860,s16861,s16862,s16863,s16864,s16865,s16866,s16867,s16868,s16869,s16870,s16871,s16872,s16873,s16874,s16875,s16876,s16877,s16878,s16879,

s16880,s16881,s16882,s16883,s16884,s16885,s16886,s16887,s16888,s16889,s16890,s16891,s16892,s16893,s16894,s16895,
	a1,b1,c1,d1,
	a2,b2,c2,d2,
	a3,b3,c3,d3,
	a4,b4,c4,d4,
	a5,b5,c5,d5,
	a6,b6,c6,d6,
	a7,b7,c7,d7,
	a8,b8,c8,d8,
	ab1,ab2,ab3,ab4,ab5,ab6,ab7,ab8,
	ab9,ab10,ab11,ab12,ab13,ab14,ab15,ab16,
	ab17,ab18,ab19,ab20,ab21,ab22,ab23,ab24,
	calculate,calculate0,
	calculate00,calculate01,calculate02,calculate03,
	calculate04,calculate05,calculate06,calculate07,
	calculate1,calculate2,calculate3,calculate4,calculate5,
	calculate6,calculate7,calculate8,calculate9,calculate10,
	calculate11,calculate12,calculate13,calculate14,calculate15,
	calculate16,calculate17,calculate18,calculate19,calculate20,
	ending0,ending1,ending2,ending);
	variable state : states;
	variable voccRemScale : std_logic_vector (31 downto 0);
	variable voccColumnScale : std_logic_vector (31 downto 0);
	variable voccRowScale : std_logic_vector (31 downto 0);

	variable voccRemScale1 : std_logic_vector (3 downto 0);
	variable voccColumnScale1 : std_logic_vector (3 downto 0);
	variable voccRowScale1 : std_logic_vector (3 downto 0);

	variable voffsetRef1: std_logic_vector (15 downto 0);
	variable voffsetRef : std_logic_vector (15 downto 0);
	variable fptmp1,fptmp2 : std_logic_vector (31 downto 0);
	variable row,col,vocccolumnj,occrowi,voccrowi,vOffsetAverage,voffset_ft : std_logic_vector (31 downto 0);
	variable temp1,voffset : std_logic_vector (15 downto 0);

	variable fracas : fracas;
	variable fracbs : fracbs;
	variable fracau : fracau;
	variable fracbu : fracbu;
	variable vOffset_sf,voffsetRef_sf : st_sfixed_max;
	variable eeprom16slv,ram16slv : slv16;
	variable eeprom16sf,ram16sf : sfixed16;
	variable eeprom16uf,ram16uf : ufixed16;
begin
	if (rising_edge (i_clock)) then
		if (i_reset = '1') then
			state := idle;
			nibble1 <= (others => '0');
			nibble2 <= (others => '0');
			nibble3 <= (others => '0');
			i := 0;
			j := 0;
			write_enable <= '0';
			ena_mux1 <= '0';
			rdy <= '0';
			addfpsclr <= '1';
			mulfpsclr <= '1';
			fixed2floatsclr <= '1';
			mulfpa <= (others => '0');
			mulfpb <= (others => '0');
			addfpa <= (others => '0');
			addfpb <= (others => '0');
			addfpond <= '0';
			mulfpond <= '0';
			addfpce <= '0';
			mulfpce <= '0';
			addra <= (others => '0');
			dia <= (others => '0');
			o_done <= '0';
			i2c_mem_ena <= '0';
		else
			case (state) is
				when idle =>
					if (i_run = '1') then
						state := occ0;
						i2c_mem_ena <= '1';
						write_enable <= '1';
						ena_mux1 <= '1';
					else
						state := idle;
						i2c_mem_ena <= '0';
						write_enable <= '0';
						ena_mux1 <= '0';
					end if;
				when occ0 => state := occ1;
					i := 0; j := 0;
					addfpsclr <= '0';
					mulfpsclr <= '0';
					fixed2floatsclr <= '0';
					rdy <= '0';
					
				when occ1 => state := occ2;
					i2c_mem_addra <= std_logic_vector (to_unsigned (0, 12)); -- 2410 LSB
				when occ2 => state := occ3;
					i2c_mem_addra <= std_logic_vector (to_unsigned (1, 12)); -- 2410 MSB
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ3 => state := occ4;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ4 => state := occ5;
					nibble1 <= temp1 (3 downto 0); -- occ scale remnant
				when occ5 => state := occ6;
				
					voccRemScale := out_nibble1; -- out occ scale remnant signed
					voccRemScale1 := temp1 (3 downto 0); -- occ scale remnant for 2^x
					
					nibble1 <= temp1 (7 downto 4); -- occ scale column
				when occ6 => state := occ7;
				
					voccColumnScale := out_nibble1; -- out occ scale column signed
					voccColumnScale1 := temp1 (7 downto 4); -- occ scale column for 2^x

					nibble1 <= temp1 (11 downto 8); -- occ scale row
				when occ7 => state := occ8;
					
					voccRowScale := out_nibble1; -- out occ row column signed
					voccRowScale1 := temp1 (11 downto 8); -- occ scale row for 2^x

				when occ8 => state := occ9;
					i2c_mem_addra <= std_logic_vector (to_unsigned (2, 12)); -- 2411 LSB
				when occ9 => state := occ10;
					i2c_mem_addra <= std_logic_vector (to_unsigned (3, 12)); -- 2411 MSB
					voffsetRef (7 downto 0) := i2c_mem_douta; -- offsetref LSB
				when occ10 => state := occ11;
					voffsetRef (15 downto 8) := i2c_mem_douta; -- offsetref MSB
				
				
					
				when occ11 => state := occ12;
					i2c_mem_addra <= std_logic_vector (to_unsigned (4, 12)); -- 2412 LSB -- occrow1-4
				when occ12 => state := occ13;
					i2c_mem_addra <= std_logic_vector (to_unsigned (5, 12)); -- 2412 MSB -- occrow1-4
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ13 => state := occ14;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ14 => state := occ15;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ15 => state := occ16;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (0, 10));
				when occ16 => state := occ17;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (1, 10));
				when occ17 => state := occ18;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (2, 10));
				when occ18 => state := occ19;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (3, 10));




				when occ19 => state := occ20;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (6, 12)); -- 2413 LSB -- occrow5-8
				when occ20 => state := occ21;
					i2c_mem_addra <= std_logic_vector (to_unsigned (7, 12)); -- 2413 MSB -- occrow5-8
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ21 => state := occ22;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ22 => state := occ23;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ23 => state := occ24;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (4, 10));
				when occ24 => state := occ25;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (5, 10));
				when occ25 => state := occ26;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (6, 10));
				when occ26 => state := occ27;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (7, 10));


				when occ27 => state := occ28;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (8, 12)); -- 2414 LSB -- occrow9-12
				when occ28 => state := occ29;
					i2c_mem_addra <= std_logic_vector (to_unsigned (9, 12)); -- 2414 MSB -- occrow9-12
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ29 => state := occ30;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ30 => state := occ31;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ31 => state := occ32;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (8, 10));
				when occ32 => state := occ33;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (9, 10));
				when occ33 => state := occ34;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (10, 10));
				when occ34 => state := occ35;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (11, 10));


				when occ35 => state := occ36;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (10, 12)); -- 2415 LSB -- occrow13-16
				when occ36 => state := occ37;
					i2c_mem_addra <= std_logic_vector (to_unsigned (11, 12)); -- 2415 MSB -- occrow13-16
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ37 => state := occ38;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ38 => state := occ39;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ39 => state := occ40;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (12, 10));
				when occ40 => state := occ41;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (13, 10));
				when occ41 => state := occ42;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (14, 10));
				when occ42 => state := occ43;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (15, 10));



				when occ43 => state := occ44;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (12, 12)); -- 2416 LSB -- occrow17-20
				when occ44 => state := occ45;
					i2c_mem_addra <= std_logic_vector (to_unsigned (13, 12)); -- 2416 MSB -- occrow17-20
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ45 => state := occ46;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ46 => state := occ47;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ47 => state := occ48;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (16, 10));
				when occ48 => state := occ49;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (17, 10));
				when occ49 => state := occ50;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (18, 10));
				when occ50 => state := occ51;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (19, 10));



				when occ51 => state := occ52;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (14, 12)); -- 2417 LSB -- occrow21-24
				when occ52 => state := occ53;
					i2c_mem_addra <= std_logic_vector (to_unsigned (15, 12)); -- 2417 MSB -- occrow21-24
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ53 => state := occ54;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ54 => state := occ55;
					nibble1 <= temp1 (3 downto 0); -- occrowA
				when occ55 => state := occ56;
					nibble1 <= temp1 (7 downto 4); -- occrowB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (20, 10));
				when occ56 => state := occ57;
					nibble1 <= temp1 (11 downto 8); -- occrowC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (21, 10));
				when occ57 => state := occ58;
					nibble1 <= temp1 (15 downto 12); -- occrowD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (22, 10));
				when occ58 => state := occ59;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (23, 10));


				when occ59 => state := occ60;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (16, 12)); -- 2418 LSB -- occcol1-4
				when occ60 => state := occ61;
					i2c_mem_addra <= std_logic_vector (to_unsigned (17, 12)); -- 2418 MSB -- occcol1-4
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ61 => state := occ62;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ62 => state := occ63;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ63 => state := occ64;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (24, 10));
				when occ64 => state := occ65;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (25, 10));
				when occ65 => state := occ66;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (26, 10));
				when occ66 => state := occ67;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (27, 10));


				when occ67 => state := occ68;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (18, 12)); -- 2419 LSB -- occcol5-8
				when occ68 => state := occ69;
					i2c_mem_addra <= std_logic_vector (to_unsigned (19, 12)); -- 2419 MSB -- occcol5-8
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ69 => state := occ70;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ70 => state := occ71;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ71 => state := occ72;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (28, 10));
				when occ72 => state := occ73;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (29, 10));
				when occ73 => state := occ74;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (30, 10));
				when occ74 => state := occ75;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (31, 10));



				when occ75 => state := occ76;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (20, 12)); -- 241a LSB -- occcol9-12
				when occ76 => state := occ77;
					i2c_mem_addra <= std_logic_vector (to_unsigned (21, 12)); -- 241a MSB -- occcol9-12
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ77 => state := occ78;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ78 => state := occ79;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ79 => state := occ80;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (32, 10));
				when occ80 => state := occ81;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (33, 10));
				when occ81 => state := occ82;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (34, 10));
				when occ82 => state := occ83;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (35, 10));




				when occ83 => state := occ84;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (22, 12)); -- 241b LSB -- occcol13-16
				when occ84 => state := occ85;
					i2c_mem_addra <= std_logic_vector (to_unsigned (23, 12)); -- 241b MSB -- occcol13-16
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ85 => state := occ86;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ86 => state := occ87;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ87 => state := occ88;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (36, 10));
				when occ88 => state := occ89;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (37, 10));
				when occ89 => state := occ90;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (38, 10));
				when occ90 => state := occ91;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (39, 10));



				when occ91 => state := occ92;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (24, 12)); -- 241c LSB -- occcol17-20
				when occ92 => state := occ93;
					i2c_mem_addra <= std_logic_vector (to_unsigned (25, 12)); -- 241c MSB -- occcol17-20
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ93 => state := occ94;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ94 => state := occ95;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ95 => state := occ96;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (40, 10));
				when occ96 => state := occ97;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (41, 10));
				when occ97 => state := occ98;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (42, 10));
				when occ98 => state := occ99;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (43, 10));



				when occ99 => state := occ100;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (26, 12)); -- 241d LSB -- occcol21-24
				when occ100 => state := occ101;
					i2c_mem_addra <= std_logic_vector (to_unsigned (27, 12)); -- 241d MSB -- occcol21-24
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ101 => state := occ102;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ102 => state := occ103;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ103 => state := occ104;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (44, 10));
				when occ104 => state := occ105;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (45, 10));
				when occ105 => state := occ106;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (46, 10));
				when occ106 => state := occ107;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (47, 10));



				when occ107 => state := occ108;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (28, 12)); -- 241e LSB -- occcol25-28
				when occ108 => state := occ109;
					i2c_mem_addra <= std_logic_vector (to_unsigned (29, 12)); -- 241e MSB -- occcol25-28
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ109 => state := occ110;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ110 => state := occ111;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ111 => state := occ112;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (48, 10));
				when occ112 => state := occ113;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (49, 10));
				when occ113 => state := occ114;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (50, 10));
				when occ114 => state := occ115;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (51, 10));



				when occ115 => state := occ116;
					addra <= (others => '0');
					i2c_mem_addra <= std_logic_vector (to_unsigned (30, 12)); -- 241f LSB -- occcol29-32
				when occ116 => state := occ117;
					i2c_mem_addra <= std_logic_vector (to_unsigned (31, 12)); -- 241f MSB -- occcol29-32
					temp1 (7 downto 0) := i2c_mem_douta;
				when occ117 => state := occ118;
					temp1 (15 downto 8) := i2c_mem_douta;
				when occ118 => state := occ119;
					nibble1 <= temp1 (3 downto 0); -- occcolA
				when occ119 => state := occ120;
					nibble1 <= temp1 (7 downto 4); -- occcolB
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (52, 10));
				when occ120 => state := occ121;
					nibble1 <= temp1 (11 downto 8); -- occcolC
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (53, 10));
				when occ121 => state := occ122;
					nibble1 <= temp1 (15 downto 12); -- occcolD
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (54, 10));
				when occ122 => state := pow0;
					dia <= out_nibble1;
					addra <= std_logic_vector (to_unsigned (55, 10));



				when pow0 => state := pow1;
					nibble4 <= voccRemScale1;
				when pow1 => state := pow2;
					voccRemScale := out_nibble4; -- 2^occscaleremnant
					nibble4 <= voccColumnScale1;
				when pow2 => state := pow3;
					voccColumnScale := out_nibble4; -- 2^occscalecolumn
					nibble4 <= voccRowScale1;
				when pow3 => state := pow4;
					voccRowScale := out_nibble4; -- 2^occscalerow
					voffsetRef_sf := resize (to_sfixed (voffsetRef, eeprom16sf), voffsetRef_sf);
					fixed2floatce <= '1';
					fixed2floatond <= '1';
					fixed2floata <= 
					to_slv (to_sfixed (to_slv (voffsetRef_sf (fracas'high downto fracas'low)), fracas))&
					to_slv (to_sfixed (to_slv (voffsetRef_sf (fracbs'high downto fracbs'low)), fracbs));
				when pow4 =>
					if (fixed2floatrdy = '1') then state := pow5;
						vOffsetAverage := fixed2floatr;
						fixed2floatce <= '0';
						fixed2floatond <= '0';
						fixed2floatsclr <= '1';
					else state := pow4; end if;
				when pow5 => state := s0;
					fixed2floatsclr <= '0';
					
when s0 => state := s1; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (48, 12)); -- offset LSB 0
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s1 => state := s2;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (49, 12)); -- offset MSB 1
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2 => state := s3; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3 => 			--4
	if (fixed2floatrdy = '1') then state := s4;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3; end if;
when s4 => state := s5; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5 => 			--6
	if (mulfprdy = '1') then state := s6;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5; end if;
when s6 => state := s7; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7 => 			--8
	if (mulfprdy = '1') then state := s8;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7; end if;
when s8 => state := s9; 	--9
	mulfpsclr <= '0';
when s9 => state := s10; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10 => 			--11
	if (mulfprdy = '1') then state := s11;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10; end if;
when s11 => state := s12; 	--12
	mulfpsclr <= '0';
when s12 => state := s13; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13 => 			--14
	if (addfprdy = '1') then state := s14;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13; end if;
when s14 => state := s15; 	--15
	addfpsclr <= '0';
when s15 => state := s16; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16 => 			--17
	if (addfprdy = '1') then state := s17;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16; end if;
when s17 => state := s18; 	--18
	addfpsclr <= '0';
when s18 => state := s19; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s19 => 			--20
	if (addfprdy = '1') then state := s20;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s19; end if;
when s20 => state := s21; 	--21
	addfpsclr <= '0';
when s21 => state := s22; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (56, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s22 => state := s23; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (50, 12)); -- offset LSB 2
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s23 => state := s24;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (51, 12)); -- offset MSB 3
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s24 => state := s25; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s25 => 			--4
	if (fixed2floatrdy = '1') then state := s26;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s25; end if;
when s26 => state := s27; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s27 => 			--6
	if (mulfprdy = '1') then state := s28;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s27; end if;
when s28 => state := s29; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s29 => 			--8
	if (mulfprdy = '1') then state := s30;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s29; end if;
when s30 => state := s31; 	--9
	mulfpsclr <= '0';
when s31 => state := s32; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s32 => 			--11
	if (mulfprdy = '1') then state := s33;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s32; end if;
when s33 => state := s34; 	--12
	mulfpsclr <= '0';
when s34 => state := s35; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s35 => 			--14
	if (addfprdy = '1') then state := s36;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s35; end if;
when s36 => state := s37; 	--15
	addfpsclr <= '0';
when s37 => state := s38; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s38 => 			--17
	if (addfprdy = '1') then state := s39;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s38; end if;
when s39 => state := s40; 	--18
	addfpsclr <= '0';
when s40 => state := s41; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s41 => 			--20
	if (addfprdy = '1') then state := s42;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s41; end if;
when s42 => state := s43; 	--21
	addfpsclr <= '0';
when s43 => state := s44; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (57, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s44 => state := s45; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (52, 12)); -- offset LSB 4
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s45 => state := s46;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (53, 12)); -- offset MSB 5
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s46 => state := s47; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s47 => 			--4
	if (fixed2floatrdy = '1') then state := s48;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s47; end if;
when s48 => state := s49; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s49 => 			--6
	if (mulfprdy = '1') then state := s50;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s49; end if;
when s50 => state := s51; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s51 => 			--8
	if (mulfprdy = '1') then state := s52;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s51; end if;
when s52 => state := s53; 	--9
	mulfpsclr <= '0';
when s53 => state := s54; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s54 => 			--11
	if (mulfprdy = '1') then state := s55;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s54; end if;
when s55 => state := s56; 	--12
	mulfpsclr <= '0';
when s56 => state := s57; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s57 => 			--14
	if (addfprdy = '1') then state := s58;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s57; end if;
when s58 => state := s59; 	--15
	addfpsclr <= '0';
when s59 => state := s60; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s60 => 			--17
	if (addfprdy = '1') then state := s61;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s60; end if;
when s61 => state := s62; 	--18
	addfpsclr <= '0';
when s62 => state := s63; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s63 => 			--20
	if (addfprdy = '1') then state := s64;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s63; end if;
when s64 => state := s65; 	--21
	addfpsclr <= '0';
when s65 => state := s66; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (58, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s66 => state := s67; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (54, 12)); -- offset LSB 6
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s67 => state := s68;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (55, 12)); -- offset MSB 7
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s68 => state := s69; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s69 => 			--4
	if (fixed2floatrdy = '1') then state := s70;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s69; end if;
when s70 => state := s71; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s71 => 			--6
	if (mulfprdy = '1') then state := s72;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s71; end if;
when s72 => state := s73; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s73 => 			--8
	if (mulfprdy = '1') then state := s74;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s73; end if;
when s74 => state := s75; 	--9
	mulfpsclr <= '0';
when s75 => state := s76; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s76 => 			--11
	if (mulfprdy = '1') then state := s77;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s76; end if;
when s77 => state := s78; 	--12
	mulfpsclr <= '0';
when s78 => state := s79; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s79 => 			--14
	if (addfprdy = '1') then state := s80;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s79; end if;
when s80 => state := s81; 	--15
	addfpsclr <= '0';
when s81 => state := s82; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s82 => 			--17
	if (addfprdy = '1') then state := s83;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s82; end if;
when s83 => state := s84; 	--18
	addfpsclr <= '0';
when s84 => state := s85; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s85 => 			--20
	if (addfprdy = '1') then state := s86;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s85; end if;
when s86 => state := s87; 	--21
	addfpsclr <= '0';
when s87 => state := s88; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (59, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s88 => state := s89; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (56, 12)); -- offset LSB 8
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s89 => state := s90;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (57, 12)); -- offset MSB 9
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s90 => state := s91; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s91 => 			--4
	if (fixed2floatrdy = '1') then state := s92;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s91; end if;
when s92 => state := s93; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s93 => 			--6
	if (mulfprdy = '1') then state := s94;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s93; end if;
when s94 => state := s95; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s95 => 			--8
	if (mulfprdy = '1') then state := s96;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s95; end if;
when s96 => state := s97; 	--9
	mulfpsclr <= '0';
when s97 => state := s98; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s98 => 			--11
	if (mulfprdy = '1') then state := s99;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s98; end if;
when s99 => state := s100; 	--12
	mulfpsclr <= '0';
when s100 => state := s101; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s101 => 			--14
	if (addfprdy = '1') then state := s102;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s101; end if;
when s102 => state := s103; 	--15
	addfpsclr <= '0';
when s103 => state := s104; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s104 => 			--17
	if (addfprdy = '1') then state := s105;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s104; end if;
when s105 => state := s106; 	--18
	addfpsclr <= '0';
when s106 => state := s107; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s107 => 			--20
	if (addfprdy = '1') then state := s108;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s107; end if;
when s108 => state := s109; 	--21
	addfpsclr <= '0';
when s109 => state := s110; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (60, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s110 => state := s111; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (58, 12)); -- offset LSB 10
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s111 => state := s112;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (59, 12)); -- offset MSB 11
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s112 => state := s113; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s113 => 			--4
	if (fixed2floatrdy = '1') then state := s114;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s113; end if;
when s114 => state := s115; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s115 => 			--6
	if (mulfprdy = '1') then state := s116;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s115; end if;
when s116 => state := s117; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s117 => 			--8
	if (mulfprdy = '1') then state := s118;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s117; end if;
when s118 => state := s119; 	--9
	mulfpsclr <= '0';
when s119 => state := s120; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s120 => 			--11
	if (mulfprdy = '1') then state := s121;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s120; end if;
when s121 => state := s122; 	--12
	mulfpsclr <= '0';
when s122 => state := s123; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s123 => 			--14
	if (addfprdy = '1') then state := s124;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s123; end if;
when s124 => state := s125; 	--15
	addfpsclr <= '0';
when s125 => state := s126; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s126 => 			--17
	if (addfprdy = '1') then state := s127;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s126; end if;
when s127 => state := s128; 	--18
	addfpsclr <= '0';
when s128 => state := s129; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s129 => 			--20
	if (addfprdy = '1') then state := s130;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s129; end if;
when s130 => state := s131; 	--21
	addfpsclr <= '0';
when s131 => state := s132; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (61, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s132 => state := s133; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (60, 12)); -- offset LSB 12
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s133 => state := s134;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (61, 12)); -- offset MSB 13
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s134 => state := s135; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s135 => 			--4
	if (fixed2floatrdy = '1') then state := s136;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s135; end if;
when s136 => state := s137; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s137 => 			--6
	if (mulfprdy = '1') then state := s138;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s137; end if;
when s138 => state := s139; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s139 => 			--8
	if (mulfprdy = '1') then state := s140;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s139; end if;
when s140 => state := s141; 	--9
	mulfpsclr <= '0';
when s141 => state := s142; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s142 => 			--11
	if (mulfprdy = '1') then state := s143;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s142; end if;
when s143 => state := s144; 	--12
	mulfpsclr <= '0';
when s144 => state := s145; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s145 => 			--14
	if (addfprdy = '1') then state := s146;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s145; end if;
when s146 => state := s147; 	--15
	addfpsclr <= '0';
when s147 => state := s148; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s148 => 			--17
	if (addfprdy = '1') then state := s149;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s148; end if;
when s149 => state := s150; 	--18
	addfpsclr <= '0';
when s150 => state := s151; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s151 => 			--20
	if (addfprdy = '1') then state := s152;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s151; end if;
when s152 => state := s153; 	--21
	addfpsclr <= '0';
when s153 => state := s154; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (62, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s154 => state := s155; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (62, 12)); -- offset LSB 14
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s155 => state := s156;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (63, 12)); -- offset MSB 15
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s156 => state := s157; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s157 => 			--4
	if (fixed2floatrdy = '1') then state := s158;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s157; end if;
when s158 => state := s159; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s159 => 			--6
	if (mulfprdy = '1') then state := s160;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s159; end if;
when s160 => state := s161; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s161 => 			--8
	if (mulfprdy = '1') then state := s162;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s161; end if;
when s162 => state := s163; 	--9
	mulfpsclr <= '0';
when s163 => state := s164; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s164 => 			--11
	if (mulfprdy = '1') then state := s165;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s164; end if;
when s165 => state := s166; 	--12
	mulfpsclr <= '0';
when s166 => state := s167; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s167 => 			--14
	if (addfprdy = '1') then state := s168;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s167; end if;
when s168 => state := s169; 	--15
	addfpsclr <= '0';
when s169 => state := s170; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s170 => 			--17
	if (addfprdy = '1') then state := s171;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s170; end if;
when s171 => state := s172; 	--18
	addfpsclr <= '0';
when s172 => state := s173; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s173 => 			--20
	if (addfprdy = '1') then state := s174;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s173; end if;
when s174 => state := s175; 	--21
	addfpsclr <= '0';
when s175 => state := s176; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (63, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s176 => state := s177; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (64, 12)); -- offset LSB 16
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s177 => state := s178;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (65, 12)); -- offset MSB 17
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s178 => state := s179; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s179 => 			--4
	if (fixed2floatrdy = '1') then state := s180;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s179; end if;
when s180 => state := s181; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s181 => 			--6
	if (mulfprdy = '1') then state := s182;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s181; end if;
when s182 => state := s183; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s183 => 			--8
	if (mulfprdy = '1') then state := s184;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s183; end if;
when s184 => state := s185; 	--9
	mulfpsclr <= '0';
when s185 => state := s186; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s186 => 			--11
	if (mulfprdy = '1') then state := s187;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s186; end if;
when s187 => state := s188; 	--12
	mulfpsclr <= '0';
when s188 => state := s189; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s189 => 			--14
	if (addfprdy = '1') then state := s190;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s189; end if;
when s190 => state := s191; 	--15
	addfpsclr <= '0';
when s191 => state := s192; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s192 => 			--17
	if (addfprdy = '1') then state := s193;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s192; end if;
when s193 => state := s194; 	--18
	addfpsclr <= '0';
when s194 => state := s195; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s195 => 			--20
	if (addfprdy = '1') then state := s196;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s195; end if;
when s196 => state := s197; 	--21
	addfpsclr <= '0';
when s197 => state := s198; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (64, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s198 => state := s199; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (66, 12)); -- offset LSB 18
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s199 => state := s200;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (67, 12)); -- offset MSB 19
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s200 => state := s201; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s201 => 			--4
	if (fixed2floatrdy = '1') then state := s202;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s201; end if;
when s202 => state := s203; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s203 => 			--6
	if (mulfprdy = '1') then state := s204;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s203; end if;
when s204 => state := s205; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s205 => 			--8
	if (mulfprdy = '1') then state := s206;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s205; end if;
when s206 => state := s207; 	--9
	mulfpsclr <= '0';
when s207 => state := s208; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s208 => 			--11
	if (mulfprdy = '1') then state := s209;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s208; end if;
when s209 => state := s210; 	--12
	mulfpsclr <= '0';
when s210 => state := s211; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s211 => 			--14
	if (addfprdy = '1') then state := s212;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s211; end if;
when s212 => state := s213; 	--15
	addfpsclr <= '0';
when s213 => state := s214; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s214 => 			--17
	if (addfprdy = '1') then state := s215;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s214; end if;
when s215 => state := s216; 	--18
	addfpsclr <= '0';
when s216 => state := s217; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s217 => 			--20
	if (addfprdy = '1') then state := s218;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s217; end if;
when s218 => state := s219; 	--21
	addfpsclr <= '0';
when s219 => state := s220; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (65, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s220 => state := s221; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (68, 12)); -- offset LSB 20
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s221 => state := s222;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (69, 12)); -- offset MSB 21
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s222 => state := s223; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s223 => 			--4
	if (fixed2floatrdy = '1') then state := s224;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s223; end if;
when s224 => state := s225; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s225 => 			--6
	if (mulfprdy = '1') then state := s226;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s225; end if;
when s226 => state := s227; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s227 => 			--8
	if (mulfprdy = '1') then state := s228;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s227; end if;
when s228 => state := s229; 	--9
	mulfpsclr <= '0';
when s229 => state := s230; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s230 => 			--11
	if (mulfprdy = '1') then state := s231;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s230; end if;
when s231 => state := s232; 	--12
	mulfpsclr <= '0';
when s232 => state := s233; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s233 => 			--14
	if (addfprdy = '1') then state := s234;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s233; end if;
when s234 => state := s235; 	--15
	addfpsclr <= '0';
when s235 => state := s236; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s236 => 			--17
	if (addfprdy = '1') then state := s237;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s236; end if;
when s237 => state := s238; 	--18
	addfpsclr <= '0';
when s238 => state := s239; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s239 => 			--20
	if (addfprdy = '1') then state := s240;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s239; end if;
when s240 => state := s241; 	--21
	addfpsclr <= '0';
when s241 => state := s242; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (66, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s242 => state := s243; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (70, 12)); -- offset LSB 22
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s243 => state := s244;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (71, 12)); -- offset MSB 23
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s244 => state := s245; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s245 => 			--4
	if (fixed2floatrdy = '1') then state := s246;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s245; end if;
when s246 => state := s247; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s247 => 			--6
	if (mulfprdy = '1') then state := s248;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s247; end if;
when s248 => state := s249; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s249 => 			--8
	if (mulfprdy = '1') then state := s250;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s249; end if;
when s250 => state := s251; 	--9
	mulfpsclr <= '0';
when s251 => state := s252; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s252 => 			--11
	if (mulfprdy = '1') then state := s253;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s252; end if;
when s253 => state := s254; 	--12
	mulfpsclr <= '0';
when s254 => state := s255; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s255 => 			--14
	if (addfprdy = '1') then state := s256;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s255; end if;
when s256 => state := s257; 	--15
	addfpsclr <= '0';
when s257 => state := s258; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s258 => 			--17
	if (addfprdy = '1') then state := s259;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s258; end if;
when s259 => state := s260; 	--18
	addfpsclr <= '0';
when s260 => state := s261; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s261 => 			--20
	if (addfprdy = '1') then state := s262;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s261; end if;
when s262 => state := s263; 	--21
	addfpsclr <= '0';
when s263 => state := s264; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (67, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s264 => state := s265; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (72, 12)); -- offset LSB 24
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s265 => state := s266;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (73, 12)); -- offset MSB 25
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s266 => state := s267; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s267 => 			--4
	if (fixed2floatrdy = '1') then state := s268;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s267; end if;
when s268 => state := s269; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s269 => 			--6
	if (mulfprdy = '1') then state := s270;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s269; end if;
when s270 => state := s271; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s271 => 			--8
	if (mulfprdy = '1') then state := s272;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s271; end if;
when s272 => state := s273; 	--9
	mulfpsclr <= '0';
when s273 => state := s274; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s274 => 			--11
	if (mulfprdy = '1') then state := s275;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s274; end if;
when s275 => state := s276; 	--12
	mulfpsclr <= '0';
when s276 => state := s277; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s277 => 			--14
	if (addfprdy = '1') then state := s278;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s277; end if;
when s278 => state := s279; 	--15
	addfpsclr <= '0';
when s279 => state := s280; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s280 => 			--17
	if (addfprdy = '1') then state := s281;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s280; end if;
when s281 => state := s282; 	--18
	addfpsclr <= '0';
when s282 => state := s283; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s283 => 			--20
	if (addfprdy = '1') then state := s284;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s283; end if;
when s284 => state := s285; 	--21
	addfpsclr <= '0';
when s285 => state := s286; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (68, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s286 => state := s287; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (74, 12)); -- offset LSB 26
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s287 => state := s288;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (75, 12)); -- offset MSB 27
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s288 => state := s289; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s289 => 			--4
	if (fixed2floatrdy = '1') then state := s290;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s289; end if;
when s290 => state := s291; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s291 => 			--6
	if (mulfprdy = '1') then state := s292;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s291; end if;
when s292 => state := s293; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s293 => 			--8
	if (mulfprdy = '1') then state := s294;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s293; end if;
when s294 => state := s295; 	--9
	mulfpsclr <= '0';
when s295 => state := s296; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s296 => 			--11
	if (mulfprdy = '1') then state := s297;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s296; end if;
when s297 => state := s298; 	--12
	mulfpsclr <= '0';
when s298 => state := s299; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s299 => 			--14
	if (addfprdy = '1') then state := s300;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s299; end if;
when s300 => state := s301; 	--15
	addfpsclr <= '0';
when s301 => state := s302; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s302 => 			--17
	if (addfprdy = '1') then state := s303;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s302; end if;
when s303 => state := s304; 	--18
	addfpsclr <= '0';
when s304 => state := s305; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s305 => 			--20
	if (addfprdy = '1') then state := s306;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s305; end if;
when s306 => state := s307; 	--21
	addfpsclr <= '0';
when s307 => state := s308; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (69, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s308 => state := s309; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (76, 12)); -- offset LSB 28
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s309 => state := s310;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (77, 12)); -- offset MSB 29
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s310 => state := s311; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s311 => 			--4
	if (fixed2floatrdy = '1') then state := s312;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s311; end if;
when s312 => state := s313; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s313 => 			--6
	if (mulfprdy = '1') then state := s314;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s313; end if;
when s314 => state := s315; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s315 => 			--8
	if (mulfprdy = '1') then state := s316;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s315; end if;
when s316 => state := s317; 	--9
	mulfpsclr <= '0';
when s317 => state := s318; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s318 => 			--11
	if (mulfprdy = '1') then state := s319;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s318; end if;
when s319 => state := s320; 	--12
	mulfpsclr <= '0';
when s320 => state := s321; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s321 => 			--14
	if (addfprdy = '1') then state := s322;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s321; end if;
when s322 => state := s323; 	--15
	addfpsclr <= '0';
when s323 => state := s324; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s324 => 			--17
	if (addfprdy = '1') then state := s325;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s324; end if;
when s325 => state := s326; 	--18
	addfpsclr <= '0';
when s326 => state := s327; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s327 => 			--20
	if (addfprdy = '1') then state := s328;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s327; end if;
when s328 => state := s329; 	--21
	addfpsclr <= '0';
when s329 => state := s330; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (70, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s330 => state := s331; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (78, 12)); -- offset LSB 30
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s331 => state := s332;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (79, 12)); -- offset MSB 31
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s332 => state := s333; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s333 => 			--4
	if (fixed2floatrdy = '1') then state := s334;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s333; end if;
when s334 => state := s335; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s335 => 			--6
	if (mulfprdy = '1') then state := s336;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s335; end if;
when s336 => state := s337; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s337 => 			--8
	if (mulfprdy = '1') then state := s338;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s337; end if;
when s338 => state := s339; 	--9
	mulfpsclr <= '0';
when s339 => state := s340; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s340 => 			--11
	if (mulfprdy = '1') then state := s341;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s340; end if;
when s341 => state := s342; 	--12
	mulfpsclr <= '0';
when s342 => state := s343; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s343 => 			--14
	if (addfprdy = '1') then state := s344;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s343; end if;
when s344 => state := s345; 	--15
	addfpsclr <= '0';
when s345 => state := s346; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s346 => 			--17
	if (addfprdy = '1') then state := s347;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s346; end if;
when s347 => state := s348; 	--18
	addfpsclr <= '0';
when s348 => state := s349; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s349 => 			--20
	if (addfprdy = '1') then state := s350;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s349; end if;
when s350 => state := s351; 	--21
	addfpsclr <= '0';
when s351 => state := s352; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (71, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s352 => state := s353; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (80, 12)); -- offset LSB 32
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s353 => state := s354;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (81, 12)); -- offset MSB 33
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s354 => state := s355; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s355 => 			--4
	if (fixed2floatrdy = '1') then state := s356;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s355; end if;
when s356 => state := s357; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s357 => 			--6
	if (mulfprdy = '1') then state := s358;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s357; end if;
when s358 => state := s359; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s359 => 			--8
	if (mulfprdy = '1') then state := s360;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s359; end if;
when s360 => state := s361; 	--9
	mulfpsclr <= '0';
when s361 => state := s362; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s362 => 			--11
	if (mulfprdy = '1') then state := s363;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s362; end if;
when s363 => state := s364; 	--12
	mulfpsclr <= '0';
when s364 => state := s365; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s365 => 			--14
	if (addfprdy = '1') then state := s366;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s365; end if;
when s366 => state := s367; 	--15
	addfpsclr <= '0';
when s367 => state := s368; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s368 => 			--17
	if (addfprdy = '1') then state := s369;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s368; end if;
when s369 => state := s370; 	--18
	addfpsclr <= '0';
when s370 => state := s371; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s371 => 			--20
	if (addfprdy = '1') then state := s372;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s371; end if;
when s372 => state := s373; 	--21
	addfpsclr <= '0';
when s373 => state := s374; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (72, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s374 => state := s375; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (82, 12)); -- offset LSB 34
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s375 => state := s376;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (83, 12)); -- offset MSB 35
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s376 => state := s377; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s377 => 			--4
	if (fixed2floatrdy = '1') then state := s378;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s377; end if;
when s378 => state := s379; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s379 => 			--6
	if (mulfprdy = '1') then state := s380;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s379; end if;
when s380 => state := s381; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s381 => 			--8
	if (mulfprdy = '1') then state := s382;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s381; end if;
when s382 => state := s383; 	--9
	mulfpsclr <= '0';
when s383 => state := s384; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s384 => 			--11
	if (mulfprdy = '1') then state := s385;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s384; end if;
when s385 => state := s386; 	--12
	mulfpsclr <= '0';
when s386 => state := s387; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s387 => 			--14
	if (addfprdy = '1') then state := s388;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s387; end if;
when s388 => state := s389; 	--15
	addfpsclr <= '0';
when s389 => state := s390; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s390 => 			--17
	if (addfprdy = '1') then state := s391;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s390; end if;
when s391 => state := s392; 	--18
	addfpsclr <= '0';
when s392 => state := s393; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s393 => 			--20
	if (addfprdy = '1') then state := s394;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s393; end if;
when s394 => state := s395; 	--21
	addfpsclr <= '0';
when s395 => state := s396; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (73, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s396 => state := s397; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (84, 12)); -- offset LSB 36
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s397 => state := s398;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (85, 12)); -- offset MSB 37
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s398 => state := s399; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s399 => 			--4
	if (fixed2floatrdy = '1') then state := s400;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s399; end if;
when s400 => state := s401; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s401 => 			--6
	if (mulfprdy = '1') then state := s402;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s401; end if;
when s402 => state := s403; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s403 => 			--8
	if (mulfprdy = '1') then state := s404;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s403; end if;
when s404 => state := s405; 	--9
	mulfpsclr <= '0';
when s405 => state := s406; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s406 => 			--11
	if (mulfprdy = '1') then state := s407;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s406; end if;
when s407 => state := s408; 	--12
	mulfpsclr <= '0';
when s408 => state := s409; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s409 => 			--14
	if (addfprdy = '1') then state := s410;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s409; end if;
when s410 => state := s411; 	--15
	addfpsclr <= '0';
when s411 => state := s412; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s412 => 			--17
	if (addfprdy = '1') then state := s413;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s412; end if;
when s413 => state := s414; 	--18
	addfpsclr <= '0';
when s414 => state := s415; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s415 => 			--20
	if (addfprdy = '1') then state := s416;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s415; end if;
when s416 => state := s417; 	--21
	addfpsclr <= '0';
when s417 => state := s418; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (74, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s418 => state := s419; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (86, 12)); -- offset LSB 38
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s419 => state := s420;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (87, 12)); -- offset MSB 39
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s420 => state := s421; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s421 => 			--4
	if (fixed2floatrdy = '1') then state := s422;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s421; end if;
when s422 => state := s423; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s423 => 			--6
	if (mulfprdy = '1') then state := s424;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s423; end if;
when s424 => state := s425; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s425 => 			--8
	if (mulfprdy = '1') then state := s426;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s425; end if;
when s426 => state := s427; 	--9
	mulfpsclr <= '0';
when s427 => state := s428; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s428 => 			--11
	if (mulfprdy = '1') then state := s429;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s428; end if;
when s429 => state := s430; 	--12
	mulfpsclr <= '0';
when s430 => state := s431; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s431 => 			--14
	if (addfprdy = '1') then state := s432;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s431; end if;
when s432 => state := s433; 	--15
	addfpsclr <= '0';
when s433 => state := s434; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s434 => 			--17
	if (addfprdy = '1') then state := s435;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s434; end if;
when s435 => state := s436; 	--18
	addfpsclr <= '0';
when s436 => state := s437; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s437 => 			--20
	if (addfprdy = '1') then state := s438;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s437; end if;
when s438 => state := s439; 	--21
	addfpsclr <= '0';
when s439 => state := s440; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (75, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s440 => state := s441; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (88, 12)); -- offset LSB 40
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s441 => state := s442;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (89, 12)); -- offset MSB 41
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s442 => state := s443; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s443 => 			--4
	if (fixed2floatrdy = '1') then state := s444;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s443; end if;
when s444 => state := s445; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s445 => 			--6
	if (mulfprdy = '1') then state := s446;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s445; end if;
when s446 => state := s447; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s447 => 			--8
	if (mulfprdy = '1') then state := s448;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s447; end if;
when s448 => state := s449; 	--9
	mulfpsclr <= '0';
when s449 => state := s450; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s450 => 			--11
	if (mulfprdy = '1') then state := s451;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s450; end if;
when s451 => state := s452; 	--12
	mulfpsclr <= '0';
when s452 => state := s453; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s453 => 			--14
	if (addfprdy = '1') then state := s454;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s453; end if;
when s454 => state := s455; 	--15
	addfpsclr <= '0';
when s455 => state := s456; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s456 => 			--17
	if (addfprdy = '1') then state := s457;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s456; end if;
when s457 => state := s458; 	--18
	addfpsclr <= '0';
when s458 => state := s459; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s459 => 			--20
	if (addfprdy = '1') then state := s460;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s459; end if;
when s460 => state := s461; 	--21
	addfpsclr <= '0';
when s461 => state := s462; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (76, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s462 => state := s463; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (90, 12)); -- offset LSB 42
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s463 => state := s464;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (91, 12)); -- offset MSB 43
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s464 => state := s465; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s465 => 			--4
	if (fixed2floatrdy = '1') then state := s466;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s465; end if;
when s466 => state := s467; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s467 => 			--6
	if (mulfprdy = '1') then state := s468;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s467; end if;
when s468 => state := s469; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s469 => 			--8
	if (mulfprdy = '1') then state := s470;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s469; end if;
when s470 => state := s471; 	--9
	mulfpsclr <= '0';
when s471 => state := s472; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s472 => 			--11
	if (mulfprdy = '1') then state := s473;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s472; end if;
when s473 => state := s474; 	--12
	mulfpsclr <= '0';
when s474 => state := s475; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s475 => 			--14
	if (addfprdy = '1') then state := s476;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s475; end if;
when s476 => state := s477; 	--15
	addfpsclr <= '0';
when s477 => state := s478; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s478 => 			--17
	if (addfprdy = '1') then state := s479;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s478; end if;
when s479 => state := s480; 	--18
	addfpsclr <= '0';
when s480 => state := s481; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s481 => 			--20
	if (addfprdy = '1') then state := s482;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s481; end if;
when s482 => state := s483; 	--21
	addfpsclr <= '0';
when s483 => state := s484; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (77, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s484 => state := s485; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (92, 12)); -- offset LSB 44
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s485 => state := s486;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (93, 12)); -- offset MSB 45
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s486 => state := s487; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s487 => 			--4
	if (fixed2floatrdy = '1') then state := s488;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s487; end if;
when s488 => state := s489; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s489 => 			--6
	if (mulfprdy = '1') then state := s490;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s489; end if;
when s490 => state := s491; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s491 => 			--8
	if (mulfprdy = '1') then state := s492;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s491; end if;
when s492 => state := s493; 	--9
	mulfpsclr <= '0';
when s493 => state := s494; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s494 => 			--11
	if (mulfprdy = '1') then state := s495;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s494; end if;
when s495 => state := s496; 	--12
	mulfpsclr <= '0';
when s496 => state := s497; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s497 => 			--14
	if (addfprdy = '1') then state := s498;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s497; end if;
when s498 => state := s499; 	--15
	addfpsclr <= '0';
when s499 => state := s500; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s500 => 			--17
	if (addfprdy = '1') then state := s501;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s500; end if;
when s501 => state := s502; 	--18
	addfpsclr <= '0';
when s502 => state := s503; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s503 => 			--20
	if (addfprdy = '1') then state := s504;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s503; end if;
when s504 => state := s505; 	--21
	addfpsclr <= '0';
when s505 => state := s506; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (78, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s506 => state := s507; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (94, 12)); -- offset LSB 46
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s507 => state := s508;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (95, 12)); -- offset MSB 47
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s508 => state := s509; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s509 => 			--4
	if (fixed2floatrdy = '1') then state := s510;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s509; end if;
when s510 => state := s511; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s511 => 			--6
	if (mulfprdy = '1') then state := s512;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s511; end if;
when s512 => state := s513; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s513 => 			--8
	if (mulfprdy = '1') then state := s514;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s513; end if;
when s514 => state := s515; 	--9
	mulfpsclr <= '0';
when s515 => state := s516; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s516 => 			--11
	if (mulfprdy = '1') then state := s517;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s516; end if;
when s517 => state := s518; 	--12
	mulfpsclr <= '0';
when s518 => state := s519; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s519 => 			--14
	if (addfprdy = '1') then state := s520;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s519; end if;
when s520 => state := s521; 	--15
	addfpsclr <= '0';
when s521 => state := s522; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s522 => 			--17
	if (addfprdy = '1') then state := s523;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s522; end if;
when s523 => state := s524; 	--18
	addfpsclr <= '0';
when s524 => state := s525; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s525 => 			--20
	if (addfprdy = '1') then state := s526;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s525; end if;
when s526 => state := s527; 	--21
	addfpsclr <= '0';
when s527 => state := s528; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (79, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s528 => state := s529; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (96, 12)); -- offset LSB 48
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s529 => state := s530;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (97, 12)); -- offset MSB 49
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s530 => state := s531; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s531 => 			--4
	if (fixed2floatrdy = '1') then state := s532;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s531; end if;
when s532 => state := s533; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s533 => 			--6
	if (mulfprdy = '1') then state := s534;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s533; end if;
when s534 => state := s535; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s535 => 			--8
	if (mulfprdy = '1') then state := s536;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s535; end if;
when s536 => state := s537; 	--9
	mulfpsclr <= '0';
when s537 => state := s538; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s538 => 			--11
	if (mulfprdy = '1') then state := s539;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s538; end if;
when s539 => state := s540; 	--12
	mulfpsclr <= '0';
when s540 => state := s541; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s541 => 			--14
	if (addfprdy = '1') then state := s542;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s541; end if;
when s542 => state := s543; 	--15
	addfpsclr <= '0';
when s543 => state := s544; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s544 => 			--17
	if (addfprdy = '1') then state := s545;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s544; end if;
when s545 => state := s546; 	--18
	addfpsclr <= '0';
when s546 => state := s547; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s547 => 			--20
	if (addfprdy = '1') then state := s548;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s547; end if;
when s548 => state := s549; 	--21
	addfpsclr <= '0';
when s549 => state := s550; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (80, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s550 => state := s551; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (98, 12)); -- offset LSB 50
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s551 => state := s552;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (99, 12)); -- offset MSB 51
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s552 => state := s553; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s553 => 			--4
	if (fixed2floatrdy = '1') then state := s554;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s553; end if;
when s554 => state := s555; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s555 => 			--6
	if (mulfprdy = '1') then state := s556;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s555; end if;
when s556 => state := s557; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s557 => 			--8
	if (mulfprdy = '1') then state := s558;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s557; end if;
when s558 => state := s559; 	--9
	mulfpsclr <= '0';
when s559 => state := s560; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s560 => 			--11
	if (mulfprdy = '1') then state := s561;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s560; end if;
when s561 => state := s562; 	--12
	mulfpsclr <= '0';
when s562 => state := s563; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s563 => 			--14
	if (addfprdy = '1') then state := s564;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s563; end if;
when s564 => state := s565; 	--15
	addfpsclr <= '0';
when s565 => state := s566; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s566 => 			--17
	if (addfprdy = '1') then state := s567;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s566; end if;
when s567 => state := s568; 	--18
	addfpsclr <= '0';
when s568 => state := s569; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s569 => 			--20
	if (addfprdy = '1') then state := s570;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s569; end if;
when s570 => state := s571; 	--21
	addfpsclr <= '0';
when s571 => state := s572; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (81, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s572 => state := s573; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (100, 12)); -- offset LSB 52
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s573 => state := s574;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (101, 12)); -- offset MSB 53
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s574 => state := s575; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s575 => 			--4
	if (fixed2floatrdy = '1') then state := s576;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s575; end if;
when s576 => state := s577; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s577 => 			--6
	if (mulfprdy = '1') then state := s578;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s577; end if;
when s578 => state := s579; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s579 => 			--8
	if (mulfprdy = '1') then state := s580;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s579; end if;
when s580 => state := s581; 	--9
	mulfpsclr <= '0';
when s581 => state := s582; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s582 => 			--11
	if (mulfprdy = '1') then state := s583;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s582; end if;
when s583 => state := s584; 	--12
	mulfpsclr <= '0';
when s584 => state := s585; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s585 => 			--14
	if (addfprdy = '1') then state := s586;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s585; end if;
when s586 => state := s587; 	--15
	addfpsclr <= '0';
when s587 => state := s588; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s588 => 			--17
	if (addfprdy = '1') then state := s589;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s588; end if;
when s589 => state := s590; 	--18
	addfpsclr <= '0';
when s590 => state := s591; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s591 => 			--20
	if (addfprdy = '1') then state := s592;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s591; end if;
when s592 => state := s593; 	--21
	addfpsclr <= '0';
when s593 => state := s594; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (82, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s594 => state := s595; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (102, 12)); -- offset LSB 54
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s595 => state := s596;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (103, 12)); -- offset MSB 55
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s596 => state := s597; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s597 => 			--4
	if (fixed2floatrdy = '1') then state := s598;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s597; end if;
when s598 => state := s599; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s599 => 			--6
	if (mulfprdy = '1') then state := s600;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s599; end if;
when s600 => state := s601; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s601 => 			--8
	if (mulfprdy = '1') then state := s602;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s601; end if;
when s602 => state := s603; 	--9
	mulfpsclr <= '0';
when s603 => state := s604; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s604 => 			--11
	if (mulfprdy = '1') then state := s605;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s604; end if;
when s605 => state := s606; 	--12
	mulfpsclr <= '0';
when s606 => state := s607; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s607 => 			--14
	if (addfprdy = '1') then state := s608;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s607; end if;
when s608 => state := s609; 	--15
	addfpsclr <= '0';
when s609 => state := s610; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s610 => 			--17
	if (addfprdy = '1') then state := s611;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s610; end if;
when s611 => state := s612; 	--18
	addfpsclr <= '0';
when s612 => state := s613; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s613 => 			--20
	if (addfprdy = '1') then state := s614;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s613; end if;
when s614 => state := s615; 	--21
	addfpsclr <= '0';
when s615 => state := s616; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (83, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s616 => state := s617; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (104, 12)); -- offset LSB 56
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s617 => state := s618;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (105, 12)); -- offset MSB 57
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s618 => state := s619; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s619 => 			--4
	if (fixed2floatrdy = '1') then state := s620;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s619; end if;
when s620 => state := s621; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s621 => 			--6
	if (mulfprdy = '1') then state := s622;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s621; end if;
when s622 => state := s623; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s623 => 			--8
	if (mulfprdy = '1') then state := s624;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s623; end if;
when s624 => state := s625; 	--9
	mulfpsclr <= '0';
when s625 => state := s626; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s626 => 			--11
	if (mulfprdy = '1') then state := s627;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s626; end if;
when s627 => state := s628; 	--12
	mulfpsclr <= '0';
when s628 => state := s629; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s629 => 			--14
	if (addfprdy = '1') then state := s630;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s629; end if;
when s630 => state := s631; 	--15
	addfpsclr <= '0';
when s631 => state := s632; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s632 => 			--17
	if (addfprdy = '1') then state := s633;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s632; end if;
when s633 => state := s634; 	--18
	addfpsclr <= '0';
when s634 => state := s635; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s635 => 			--20
	if (addfprdy = '1') then state := s636;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s635; end if;
when s636 => state := s637; 	--21
	addfpsclr <= '0';
when s637 => state := s638; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (84, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s638 => state := s639; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (106, 12)); -- offset LSB 58
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s639 => state := s640;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (107, 12)); -- offset MSB 59
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s640 => state := s641; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s641 => 			--4
	if (fixed2floatrdy = '1') then state := s642;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s641; end if;
when s642 => state := s643; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s643 => 			--6
	if (mulfprdy = '1') then state := s644;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s643; end if;
when s644 => state := s645; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s645 => 			--8
	if (mulfprdy = '1') then state := s646;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s645; end if;
when s646 => state := s647; 	--9
	mulfpsclr <= '0';
when s647 => state := s648; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s648 => 			--11
	if (mulfprdy = '1') then state := s649;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s648; end if;
when s649 => state := s650; 	--12
	mulfpsclr <= '0';
when s650 => state := s651; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s651 => 			--14
	if (addfprdy = '1') then state := s652;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s651; end if;
when s652 => state := s653; 	--15
	addfpsclr <= '0';
when s653 => state := s654; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s654 => 			--17
	if (addfprdy = '1') then state := s655;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s654; end if;
when s655 => state := s656; 	--18
	addfpsclr <= '0';
when s656 => state := s657; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s657 => 			--20
	if (addfprdy = '1') then state := s658;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s657; end if;
when s658 => state := s659; 	--21
	addfpsclr <= '0';
when s659 => state := s660; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (85, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s660 => state := s661; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (108, 12)); -- offset LSB 60
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s661 => state := s662;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (109, 12)); -- offset MSB 61
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s662 => state := s663; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s663 => 			--4
	if (fixed2floatrdy = '1') then state := s664;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s663; end if;
when s664 => state := s665; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s665 => 			--6
	if (mulfprdy = '1') then state := s666;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s665; end if;
when s666 => state := s667; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s667 => 			--8
	if (mulfprdy = '1') then state := s668;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s667; end if;
when s668 => state := s669; 	--9
	mulfpsclr <= '0';
when s669 => state := s670; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s670 => 			--11
	if (mulfprdy = '1') then state := s671;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s670; end if;
when s671 => state := s672; 	--12
	mulfpsclr <= '0';
when s672 => state := s673; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s673 => 			--14
	if (addfprdy = '1') then state := s674;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s673; end if;
when s674 => state := s675; 	--15
	addfpsclr <= '0';
when s675 => state := s676; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s676 => 			--17
	if (addfprdy = '1') then state := s677;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s676; end if;
when s677 => state := s678; 	--18
	addfpsclr <= '0';
when s678 => state := s679; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s679 => 			--20
	if (addfprdy = '1') then state := s680;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s679; end if;
when s680 => state := s681; 	--21
	addfpsclr <= '0';
when s681 => state := s682; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (86, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s682 => state := s683; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (110, 12)); -- offset LSB 62
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s683 => state := s684;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (111, 12)); -- offset MSB 63
	addra <= std_logic_vector (to_unsigned (0, 10)); -- OCCrowI 0
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s684 => state := s685; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s685 => 			--4
	if (fixed2floatrdy = '1') then state := s686;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s685; end if;
when s686 => state := s687; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s687 => 			--6
	if (mulfprdy = '1') then state := s688;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s687; end if;
when s688 => state := s689; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s689 => 			--8
	if (mulfprdy = '1') then state := s690;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s689; end if;
when s690 => state := s691; 	--9
	mulfpsclr <= '0';
when s691 => state := s692; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s692 => 			--11
	if (mulfprdy = '1') then state := s693;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s692; end if;
when s693 => state := s694; 	--12
	mulfpsclr <= '0';
when s694 => state := s695; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s695 => 			--14
	if (addfprdy = '1') then state := s696;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s695; end if;
when s696 => state := s697; 	--15
	addfpsclr <= '0';
when s697 => state := s698; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s698 => 			--17
	if (addfprdy = '1') then state := s699;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s698; end if;
when s699 => state := s700; 	--18
	addfpsclr <= '0';
when s700 => state := s701; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s701 => 			--20
	if (addfprdy = '1') then state := s702;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s701; end if;
when s702 => state := s703; 	--21
	addfpsclr <= '0';
when s703 => state := s704; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (87, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s704 => state := s705; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (112, 12)); -- offset LSB 64
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s705 => state := s706;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (113, 12)); -- offset MSB 65
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s706 => state := s707; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s707 => 			--4
	if (fixed2floatrdy = '1') then state := s708;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s707; end if;
when s708 => state := s709; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s709 => 			--6
	if (mulfprdy = '1') then state := s710;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s709; end if;
when s710 => state := s711; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s711 => 			--8
	if (mulfprdy = '1') then state := s712;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s711; end if;
when s712 => state := s713; 	--9
	mulfpsclr <= '0';
when s713 => state := s714; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s714 => 			--11
	if (mulfprdy = '1') then state := s715;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s714; end if;
when s715 => state := s716; 	--12
	mulfpsclr <= '0';
when s716 => state := s717; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s717 => 			--14
	if (addfprdy = '1') then state := s718;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s717; end if;
when s718 => state := s719; 	--15
	addfpsclr <= '0';
when s719 => state := s720; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s720 => 			--17
	if (addfprdy = '1') then state := s721;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s720; end if;
when s721 => state := s722; 	--18
	addfpsclr <= '0';
when s722 => state := s723; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s723 => 			--20
	if (addfprdy = '1') then state := s724;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s723; end if;
when s724 => state := s725; 	--21
	addfpsclr <= '0';
when s725 => state := s726; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (88, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s726 => state := s727; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (114, 12)); -- offset LSB 66
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s727 => state := s728;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (115, 12)); -- offset MSB 67
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s728 => state := s729; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s729 => 			--4
	if (fixed2floatrdy = '1') then state := s730;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s729; end if;
when s730 => state := s731; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s731 => 			--6
	if (mulfprdy = '1') then state := s732;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s731; end if;
when s732 => state := s733; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s733 => 			--8
	if (mulfprdy = '1') then state := s734;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s733; end if;
when s734 => state := s735; 	--9
	mulfpsclr <= '0';
when s735 => state := s736; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s736 => 			--11
	if (mulfprdy = '1') then state := s737;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s736; end if;
when s737 => state := s738; 	--12
	mulfpsclr <= '0';
when s738 => state := s739; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s739 => 			--14
	if (addfprdy = '1') then state := s740;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s739; end if;
when s740 => state := s741; 	--15
	addfpsclr <= '0';
when s741 => state := s742; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s742 => 			--17
	if (addfprdy = '1') then state := s743;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s742; end if;
when s743 => state := s744; 	--18
	addfpsclr <= '0';
when s744 => state := s745; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s745 => 			--20
	if (addfprdy = '1') then state := s746;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s745; end if;
when s746 => state := s747; 	--21
	addfpsclr <= '0';
when s747 => state := s748; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (89, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s748 => state := s749; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (116, 12)); -- offset LSB 68
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s749 => state := s750;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (117, 12)); -- offset MSB 69
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s750 => state := s751; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s751 => 			--4
	if (fixed2floatrdy = '1') then state := s752;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s751; end if;
when s752 => state := s753; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s753 => 			--6
	if (mulfprdy = '1') then state := s754;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s753; end if;
when s754 => state := s755; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s755 => 			--8
	if (mulfprdy = '1') then state := s756;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s755; end if;
when s756 => state := s757; 	--9
	mulfpsclr <= '0';
when s757 => state := s758; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s758 => 			--11
	if (mulfprdy = '1') then state := s759;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s758; end if;
when s759 => state := s760; 	--12
	mulfpsclr <= '0';
when s760 => state := s761; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s761 => 			--14
	if (addfprdy = '1') then state := s762;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s761; end if;
when s762 => state := s763; 	--15
	addfpsclr <= '0';
when s763 => state := s764; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s764 => 			--17
	if (addfprdy = '1') then state := s765;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s764; end if;
when s765 => state := s766; 	--18
	addfpsclr <= '0';
when s766 => state := s767; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s767 => 			--20
	if (addfprdy = '1') then state := s768;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s767; end if;
when s768 => state := s769; 	--21
	addfpsclr <= '0';
when s769 => state := s770; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (90, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s770 => state := s771; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (118, 12)); -- offset LSB 70
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s771 => state := s772;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (119, 12)); -- offset MSB 71
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s772 => state := s773; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s773 => 			--4
	if (fixed2floatrdy = '1') then state := s774;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s773; end if;
when s774 => state := s775; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s775 => 			--6
	if (mulfprdy = '1') then state := s776;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s775; end if;
when s776 => state := s777; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s777 => 			--8
	if (mulfprdy = '1') then state := s778;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s777; end if;
when s778 => state := s779; 	--9
	mulfpsclr <= '0';
when s779 => state := s780; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s780 => 			--11
	if (mulfprdy = '1') then state := s781;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s780; end if;
when s781 => state := s782; 	--12
	mulfpsclr <= '0';
when s782 => state := s783; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s783 => 			--14
	if (addfprdy = '1') then state := s784;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s783; end if;
when s784 => state := s785; 	--15
	addfpsclr <= '0';
when s785 => state := s786; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s786 => 			--17
	if (addfprdy = '1') then state := s787;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s786; end if;
when s787 => state := s788; 	--18
	addfpsclr <= '0';
when s788 => state := s789; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s789 => 			--20
	if (addfprdy = '1') then state := s790;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s789; end if;
when s790 => state := s791; 	--21
	addfpsclr <= '0';
when s791 => state := s792; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (91, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s792 => state := s793; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (120, 12)); -- offset LSB 72
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s793 => state := s794;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (121, 12)); -- offset MSB 73
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s794 => state := s795; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s795 => 			--4
	if (fixed2floatrdy = '1') then state := s796;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s795; end if;
when s796 => state := s797; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s797 => 			--6
	if (mulfprdy = '1') then state := s798;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s797; end if;
when s798 => state := s799; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s799 => 			--8
	if (mulfprdy = '1') then state := s800;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s799; end if;
when s800 => state := s801; 	--9
	mulfpsclr <= '0';
when s801 => state := s802; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s802 => 			--11
	if (mulfprdy = '1') then state := s803;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s802; end if;
when s803 => state := s804; 	--12
	mulfpsclr <= '0';
when s804 => state := s805; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s805 => 			--14
	if (addfprdy = '1') then state := s806;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s805; end if;
when s806 => state := s807; 	--15
	addfpsclr <= '0';
when s807 => state := s808; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s808 => 			--17
	if (addfprdy = '1') then state := s809;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s808; end if;
when s809 => state := s810; 	--18
	addfpsclr <= '0';
when s810 => state := s811; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s811 => 			--20
	if (addfprdy = '1') then state := s812;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s811; end if;
when s812 => state := s813; 	--21
	addfpsclr <= '0';
when s813 => state := s814; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (92, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s814 => state := s815; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (122, 12)); -- offset LSB 74
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s815 => state := s816;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (123, 12)); -- offset MSB 75
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s816 => state := s817; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s817 => 			--4
	if (fixed2floatrdy = '1') then state := s818;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s817; end if;
when s818 => state := s819; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s819 => 			--6
	if (mulfprdy = '1') then state := s820;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s819; end if;
when s820 => state := s821; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s821 => 			--8
	if (mulfprdy = '1') then state := s822;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s821; end if;
when s822 => state := s823; 	--9
	mulfpsclr <= '0';
when s823 => state := s824; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s824 => 			--11
	if (mulfprdy = '1') then state := s825;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s824; end if;
when s825 => state := s826; 	--12
	mulfpsclr <= '0';
when s826 => state := s827; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s827 => 			--14
	if (addfprdy = '1') then state := s828;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s827; end if;
when s828 => state := s829; 	--15
	addfpsclr <= '0';
when s829 => state := s830; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s830 => 			--17
	if (addfprdy = '1') then state := s831;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s830; end if;
when s831 => state := s832; 	--18
	addfpsclr <= '0';
when s832 => state := s833; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s833 => 			--20
	if (addfprdy = '1') then state := s834;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s833; end if;
when s834 => state := s835; 	--21
	addfpsclr <= '0';
when s835 => state := s836; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (93, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s836 => state := s837; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (124, 12)); -- offset LSB 76
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s837 => state := s838;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (125, 12)); -- offset MSB 77
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s838 => state := s839; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s839 => 			--4
	if (fixed2floatrdy = '1') then state := s840;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s839; end if;
when s840 => state := s841; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s841 => 			--6
	if (mulfprdy = '1') then state := s842;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s841; end if;
when s842 => state := s843; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s843 => 			--8
	if (mulfprdy = '1') then state := s844;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s843; end if;
when s844 => state := s845; 	--9
	mulfpsclr <= '0';
when s845 => state := s846; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s846 => 			--11
	if (mulfprdy = '1') then state := s847;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s846; end if;
when s847 => state := s848; 	--12
	mulfpsclr <= '0';
when s848 => state := s849; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s849 => 			--14
	if (addfprdy = '1') then state := s850;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s849; end if;
when s850 => state := s851; 	--15
	addfpsclr <= '0';
when s851 => state := s852; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s852 => 			--17
	if (addfprdy = '1') then state := s853;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s852; end if;
when s853 => state := s854; 	--18
	addfpsclr <= '0';
when s854 => state := s855; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s855 => 			--20
	if (addfprdy = '1') then state := s856;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s855; end if;
when s856 => state := s857; 	--21
	addfpsclr <= '0';
when s857 => state := s858; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (94, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s858 => state := s859; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (126, 12)); -- offset LSB 78
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s859 => state := s860;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (127, 12)); -- offset MSB 79
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s860 => state := s861; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s861 => 			--4
	if (fixed2floatrdy = '1') then state := s862;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s861; end if;
when s862 => state := s863; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s863 => 			--6
	if (mulfprdy = '1') then state := s864;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s863; end if;
when s864 => state := s865; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s865 => 			--8
	if (mulfprdy = '1') then state := s866;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s865; end if;
when s866 => state := s867; 	--9
	mulfpsclr <= '0';
when s867 => state := s868; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s868 => 			--11
	if (mulfprdy = '1') then state := s869;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s868; end if;
when s869 => state := s870; 	--12
	mulfpsclr <= '0';
when s870 => state := s871; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s871 => 			--14
	if (addfprdy = '1') then state := s872;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s871; end if;
when s872 => state := s873; 	--15
	addfpsclr <= '0';
when s873 => state := s874; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s874 => 			--17
	if (addfprdy = '1') then state := s875;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s874; end if;
when s875 => state := s876; 	--18
	addfpsclr <= '0';
when s876 => state := s877; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s877 => 			--20
	if (addfprdy = '1') then state := s878;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s877; end if;
when s878 => state := s879; 	--21
	addfpsclr <= '0';
when s879 => state := s880; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (95, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s880 => state := s881; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (128, 12)); -- offset LSB 80
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s881 => state := s882;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (129, 12)); -- offset MSB 81
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s882 => state := s883; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s883 => 			--4
	if (fixed2floatrdy = '1') then state := s884;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s883; end if;
when s884 => state := s885; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s885 => 			--6
	if (mulfprdy = '1') then state := s886;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s885; end if;
when s886 => state := s887; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s887 => 			--8
	if (mulfprdy = '1') then state := s888;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s887; end if;
when s888 => state := s889; 	--9
	mulfpsclr <= '0';
when s889 => state := s890; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s890 => 			--11
	if (mulfprdy = '1') then state := s891;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s890; end if;
when s891 => state := s892; 	--12
	mulfpsclr <= '0';
when s892 => state := s893; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s893 => 			--14
	if (addfprdy = '1') then state := s894;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s893; end if;
when s894 => state := s895; 	--15
	addfpsclr <= '0';
when s895 => state := s896; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s896 => 			--17
	if (addfprdy = '1') then state := s897;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s896; end if;
when s897 => state := s898; 	--18
	addfpsclr <= '0';
when s898 => state := s899; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s899 => 			--20
	if (addfprdy = '1') then state := s900;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s899; end if;
when s900 => state := s901; 	--21
	addfpsclr <= '0';
when s901 => state := s902; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (96, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s902 => state := s903; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (130, 12)); -- offset LSB 82
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s903 => state := s904;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (131, 12)); -- offset MSB 83
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s904 => state := s905; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s905 => 			--4
	if (fixed2floatrdy = '1') then state := s906;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s905; end if;
when s906 => state := s907; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s907 => 			--6
	if (mulfprdy = '1') then state := s908;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s907; end if;
when s908 => state := s909; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s909 => 			--8
	if (mulfprdy = '1') then state := s910;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s909; end if;
when s910 => state := s911; 	--9
	mulfpsclr <= '0';
when s911 => state := s912; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s912 => 			--11
	if (mulfprdy = '1') then state := s913;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s912; end if;
when s913 => state := s914; 	--12
	mulfpsclr <= '0';
when s914 => state := s915; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s915 => 			--14
	if (addfprdy = '1') then state := s916;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s915; end if;
when s916 => state := s917; 	--15
	addfpsclr <= '0';
when s917 => state := s918; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s918 => 			--17
	if (addfprdy = '1') then state := s919;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s918; end if;
when s919 => state := s920; 	--18
	addfpsclr <= '0';
when s920 => state := s921; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s921 => 			--20
	if (addfprdy = '1') then state := s922;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s921; end if;
when s922 => state := s923; 	--21
	addfpsclr <= '0';
when s923 => state := s924; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (97, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s924 => state := s925; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (132, 12)); -- offset LSB 84
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s925 => state := s926;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (133, 12)); -- offset MSB 85
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s926 => state := s927; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s927 => 			--4
	if (fixed2floatrdy = '1') then state := s928;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s927; end if;
when s928 => state := s929; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s929 => 			--6
	if (mulfprdy = '1') then state := s930;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s929; end if;
when s930 => state := s931; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s931 => 			--8
	if (mulfprdy = '1') then state := s932;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s931; end if;
when s932 => state := s933; 	--9
	mulfpsclr <= '0';
when s933 => state := s934; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s934 => 			--11
	if (mulfprdy = '1') then state := s935;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s934; end if;
when s935 => state := s936; 	--12
	mulfpsclr <= '0';
when s936 => state := s937; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s937 => 			--14
	if (addfprdy = '1') then state := s938;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s937; end if;
when s938 => state := s939; 	--15
	addfpsclr <= '0';
when s939 => state := s940; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s940 => 			--17
	if (addfprdy = '1') then state := s941;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s940; end if;
when s941 => state := s942; 	--18
	addfpsclr <= '0';
when s942 => state := s943; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s943 => 			--20
	if (addfprdy = '1') then state := s944;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s943; end if;
when s944 => state := s945; 	--21
	addfpsclr <= '0';
when s945 => state := s946; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (98, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s946 => state := s947; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (134, 12)); -- offset LSB 86
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s947 => state := s948;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (135, 12)); -- offset MSB 87
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s948 => state := s949; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s949 => 			--4
	if (fixed2floatrdy = '1') then state := s950;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s949; end if;
when s950 => state := s951; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s951 => 			--6
	if (mulfprdy = '1') then state := s952;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s951; end if;
when s952 => state := s953; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s953 => 			--8
	if (mulfprdy = '1') then state := s954;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s953; end if;
when s954 => state := s955; 	--9
	mulfpsclr <= '0';
when s955 => state := s956; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s956 => 			--11
	if (mulfprdy = '1') then state := s957;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s956; end if;
when s957 => state := s958; 	--12
	mulfpsclr <= '0';
when s958 => state := s959; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s959 => 			--14
	if (addfprdy = '1') then state := s960;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s959; end if;
when s960 => state := s961; 	--15
	addfpsclr <= '0';
when s961 => state := s962; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s962 => 			--17
	if (addfprdy = '1') then state := s963;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s962; end if;
when s963 => state := s964; 	--18
	addfpsclr <= '0';
when s964 => state := s965; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s965 => 			--20
	if (addfprdy = '1') then state := s966;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s965; end if;
when s966 => state := s967; 	--21
	addfpsclr <= '0';
when s967 => state := s968; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (99, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s968 => state := s969; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (136, 12)); -- offset LSB 88
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s969 => state := s970;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (137, 12)); -- offset MSB 89
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s970 => state := s971; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s971 => 			--4
	if (fixed2floatrdy = '1') then state := s972;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s971; end if;
when s972 => state := s973; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s973 => 			--6
	if (mulfprdy = '1') then state := s974;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s973; end if;
when s974 => state := s975; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s975 => 			--8
	if (mulfprdy = '1') then state := s976;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s975; end if;
when s976 => state := s977; 	--9
	mulfpsclr <= '0';
when s977 => state := s978; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s978 => 			--11
	if (mulfprdy = '1') then state := s979;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s978; end if;
when s979 => state := s980; 	--12
	mulfpsclr <= '0';
when s980 => state := s981; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s981 => 			--14
	if (addfprdy = '1') then state := s982;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s981; end if;
when s982 => state := s983; 	--15
	addfpsclr <= '0';
when s983 => state := s984; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s984 => 			--17
	if (addfprdy = '1') then state := s985;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s984; end if;
when s985 => state := s986; 	--18
	addfpsclr <= '0';
when s986 => state := s987; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s987 => 			--20
	if (addfprdy = '1') then state := s988;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s987; end if;
when s988 => state := s989; 	--21
	addfpsclr <= '0';
when s989 => state := s990; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (100, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s990 => state := s991; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (138, 12)); -- offset LSB 90
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s991 => state := s992;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (139, 12)); -- offset MSB 91
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s992 => state := s993; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s993 => 			--4
	if (fixed2floatrdy = '1') then state := s994;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s993; end if;
when s994 => state := s995; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s995 => 			--6
	if (mulfprdy = '1') then state := s996;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s995; end if;
when s996 => state := s997; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s997 => 			--8
	if (mulfprdy = '1') then state := s998;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s997; end if;
when s998 => state := s999; 	--9
	mulfpsclr <= '0';
when s999 => state := s1000; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1000 => 			--11
	if (mulfprdy = '1') then state := s1001;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1000; end if;
when s1001 => state := s1002; 	--12
	mulfpsclr <= '0';
when s1002 => state := s1003; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1003 => 			--14
	if (addfprdy = '1') then state := s1004;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1003; end if;
when s1004 => state := s1005; 	--15
	addfpsclr <= '0';
when s1005 => state := s1006; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1006 => 			--17
	if (addfprdy = '1') then state := s1007;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1006; end if;
when s1007 => state := s1008; 	--18
	addfpsclr <= '0';
when s1008 => state := s1009; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1009 => 			--20
	if (addfprdy = '1') then state := s1010;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1009; end if;
when s1010 => state := s1011; 	--21
	addfpsclr <= '0';
when s1011 => state := s1012; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (101, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1012 => state := s1013; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (140, 12)); -- offset LSB 92
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s1013 => state := s1014;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (141, 12)); -- offset MSB 93
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1014 => state := s1015; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1015 => 			--4
	if (fixed2floatrdy = '1') then state := s1016;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1015; end if;
when s1016 => state := s1017; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1017 => 			--6
	if (mulfprdy = '1') then state := s1018;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1017; end if;
when s1018 => state := s1019; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1019 => 			--8
	if (mulfprdy = '1') then state := s1020;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1019; end if;
when s1020 => state := s1021; 	--9
	mulfpsclr <= '0';
when s1021 => state := s1022; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1022 => 			--11
	if (mulfprdy = '1') then state := s1023;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1022; end if;
when s1023 => state := s1024; 	--12
	mulfpsclr <= '0';
when s1024 => state := s1025; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1025 => 			--14
	if (addfprdy = '1') then state := s1026;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1025; end if;
when s1026 => state := s1027; 	--15
	addfpsclr <= '0';
when s1027 => state := s1028; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1028 => 			--17
	if (addfprdy = '1') then state := s1029;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1028; end if;
when s1029 => state := s1030; 	--18
	addfpsclr <= '0';
when s1030 => state := s1031; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1031 => 			--20
	if (addfprdy = '1') then state := s1032;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1031; end if;
when s1032 => state := s1033; 	--21
	addfpsclr <= '0';
when s1033 => state := s1034; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (102, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1034 => state := s1035; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (142, 12)); -- offset LSB 94
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s1035 => state := s1036;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (143, 12)); -- offset MSB 95
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1036 => state := s1037; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1037 => 			--4
	if (fixed2floatrdy = '1') then state := s1038;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1037; end if;
when s1038 => state := s1039; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1039 => 			--6
	if (mulfprdy = '1') then state := s1040;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1039; end if;
when s1040 => state := s1041; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1041 => 			--8
	if (mulfprdy = '1') then state := s1042;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1041; end if;
when s1042 => state := s1043; 	--9
	mulfpsclr <= '0';
when s1043 => state := s1044; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1044 => 			--11
	if (mulfprdy = '1') then state := s1045;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1044; end if;
when s1045 => state := s1046; 	--12
	mulfpsclr <= '0';
when s1046 => state := s1047; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1047 => 			--14
	if (addfprdy = '1') then state := s1048;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1047; end if;
when s1048 => state := s1049; 	--15
	addfpsclr <= '0';
when s1049 => state := s1050; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1050 => 			--17
	if (addfprdy = '1') then state := s1051;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1050; end if;
when s1051 => state := s1052; 	--18
	addfpsclr <= '0';
when s1052 => state := s1053; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1053 => 			--20
	if (addfprdy = '1') then state := s1054;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1053; end if;
when s1054 => state := s1055; 	--21
	addfpsclr <= '0';
when s1055 => state := s1056; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (103, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1056 => state := s1057; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (144, 12)); -- offset LSB 96
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s1057 => state := s1058;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (145, 12)); -- offset MSB 97
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1058 => state := s1059; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1059 => 			--4
	if (fixed2floatrdy = '1') then state := s1060;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1059; end if;
when s1060 => state := s1061; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1061 => 			--6
	if (mulfprdy = '1') then state := s1062;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1061; end if;
when s1062 => state := s1063; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1063 => 			--8
	if (mulfprdy = '1') then state := s1064;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1063; end if;
when s1064 => state := s1065; 	--9
	mulfpsclr <= '0';
when s1065 => state := s1066; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1066 => 			--11
	if (mulfprdy = '1') then state := s1067;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1066; end if;
when s1067 => state := s1068; 	--12
	mulfpsclr <= '0';
when s1068 => state := s1069; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1069 => 			--14
	if (addfprdy = '1') then state := s1070;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1069; end if;
when s1070 => state := s1071; 	--15
	addfpsclr <= '0';
when s1071 => state := s1072; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1072 => 			--17
	if (addfprdy = '1') then state := s1073;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1072; end if;
when s1073 => state := s1074; 	--18
	addfpsclr <= '0';
when s1074 => state := s1075; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1075 => 			--20
	if (addfprdy = '1') then state := s1076;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1075; end if;
when s1076 => state := s1077; 	--21
	addfpsclr <= '0';
when s1077 => state := s1078; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (104, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1078 => state := s1079; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (146, 12)); -- offset LSB 98
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s1079 => state := s1080;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (147, 12)); -- offset MSB 99
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1080 => state := s1081; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1081 => 			--4
	if (fixed2floatrdy = '1') then state := s1082;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1081; end if;
when s1082 => state := s1083; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1083 => 			--6
	if (mulfprdy = '1') then state := s1084;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1083; end if;
when s1084 => state := s1085; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1085 => 			--8
	if (mulfprdy = '1') then state := s1086;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1085; end if;
when s1086 => state := s1087; 	--9
	mulfpsclr <= '0';
when s1087 => state := s1088; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1088 => 			--11
	if (mulfprdy = '1') then state := s1089;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1088; end if;
when s1089 => state := s1090; 	--12
	mulfpsclr <= '0';
when s1090 => state := s1091; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1091 => 			--14
	if (addfprdy = '1') then state := s1092;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1091; end if;
when s1092 => state := s1093; 	--15
	addfpsclr <= '0';
when s1093 => state := s1094; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1094 => 			--17
	if (addfprdy = '1') then state := s1095;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1094; end if;
when s1095 => state := s1096; 	--18
	addfpsclr <= '0';
when s1096 => state := s1097; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1097 => 			--20
	if (addfprdy = '1') then state := s1098;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1097; end if;
when s1098 => state := s1099; 	--21
	addfpsclr <= '0';
when s1099 => state := s1100; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (105, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1100 => state := s1101; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (148, 12)); -- offset LSB 100
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s1101 => state := s1102;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (149, 12)); -- offset MSB 101
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1102 => state := s1103; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1103 => 			--4
	if (fixed2floatrdy = '1') then state := s1104;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1103; end if;
when s1104 => state := s1105; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1105 => 			--6
	if (mulfprdy = '1') then state := s1106;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1105; end if;
when s1106 => state := s1107; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1107 => 			--8
	if (mulfprdy = '1') then state := s1108;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1107; end if;
when s1108 => state := s1109; 	--9
	mulfpsclr <= '0';
when s1109 => state := s1110; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1110 => 			--11
	if (mulfprdy = '1') then state := s1111;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1110; end if;
when s1111 => state := s1112; 	--12
	mulfpsclr <= '0';
when s1112 => state := s1113; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1113 => 			--14
	if (addfprdy = '1') then state := s1114;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1113; end if;
when s1114 => state := s1115; 	--15
	addfpsclr <= '0';
when s1115 => state := s1116; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1116 => 			--17
	if (addfprdy = '1') then state := s1117;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1116; end if;
when s1117 => state := s1118; 	--18
	addfpsclr <= '0';
when s1118 => state := s1119; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1119 => 			--20
	if (addfprdy = '1') then state := s1120;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1119; end if;
when s1120 => state := s1121; 	--21
	addfpsclr <= '0';
when s1121 => state := s1122; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (106, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1122 => state := s1123; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (150, 12)); -- offset LSB 102
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s1123 => state := s1124;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (151, 12)); -- offset MSB 103
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1124 => state := s1125; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1125 => 			--4
	if (fixed2floatrdy = '1') then state := s1126;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1125; end if;
when s1126 => state := s1127; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1127 => 			--6
	if (mulfprdy = '1') then state := s1128;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1127; end if;
when s1128 => state := s1129; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1129 => 			--8
	if (mulfprdy = '1') then state := s1130;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1129; end if;
when s1130 => state := s1131; 	--9
	mulfpsclr <= '0';
when s1131 => state := s1132; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1132 => 			--11
	if (mulfprdy = '1') then state := s1133;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1132; end if;
when s1133 => state := s1134; 	--12
	mulfpsclr <= '0';
when s1134 => state := s1135; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1135 => 			--14
	if (addfprdy = '1') then state := s1136;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1135; end if;
when s1136 => state := s1137; 	--15
	addfpsclr <= '0';
when s1137 => state := s1138; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1138 => 			--17
	if (addfprdy = '1') then state := s1139;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1138; end if;
when s1139 => state := s1140; 	--18
	addfpsclr <= '0';
when s1140 => state := s1141; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1141 => 			--20
	if (addfprdy = '1') then state := s1142;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1141; end if;
when s1142 => state := s1143; 	--21
	addfpsclr <= '0';
when s1143 => state := s1144; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (107, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1144 => state := s1145; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (152, 12)); -- offset LSB 104
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s1145 => state := s1146;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (153, 12)); -- offset MSB 105
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1146 => state := s1147; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1147 => 			--4
	if (fixed2floatrdy = '1') then state := s1148;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1147; end if;
when s1148 => state := s1149; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1149 => 			--6
	if (mulfprdy = '1') then state := s1150;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1149; end if;
when s1150 => state := s1151; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1151 => 			--8
	if (mulfprdy = '1') then state := s1152;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1151; end if;
when s1152 => state := s1153; 	--9
	mulfpsclr <= '0';
when s1153 => state := s1154; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1154 => 			--11
	if (mulfprdy = '1') then state := s1155;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1154; end if;
when s1155 => state := s1156; 	--12
	mulfpsclr <= '0';
when s1156 => state := s1157; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1157 => 			--14
	if (addfprdy = '1') then state := s1158;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1157; end if;
when s1158 => state := s1159; 	--15
	addfpsclr <= '0';
when s1159 => state := s1160; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1160 => 			--17
	if (addfprdy = '1') then state := s1161;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1160; end if;
when s1161 => state := s1162; 	--18
	addfpsclr <= '0';
when s1162 => state := s1163; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1163 => 			--20
	if (addfprdy = '1') then state := s1164;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1163; end if;
when s1164 => state := s1165; 	--21
	addfpsclr <= '0';
when s1165 => state := s1166; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (108, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1166 => state := s1167; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (154, 12)); -- offset LSB 106
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s1167 => state := s1168;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (155, 12)); -- offset MSB 107
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1168 => state := s1169; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1169 => 			--4
	if (fixed2floatrdy = '1') then state := s1170;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1169; end if;
when s1170 => state := s1171; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1171 => 			--6
	if (mulfprdy = '1') then state := s1172;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1171; end if;
when s1172 => state := s1173; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1173 => 			--8
	if (mulfprdy = '1') then state := s1174;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1173; end if;
when s1174 => state := s1175; 	--9
	mulfpsclr <= '0';
when s1175 => state := s1176; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1176 => 			--11
	if (mulfprdy = '1') then state := s1177;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1176; end if;
when s1177 => state := s1178; 	--12
	mulfpsclr <= '0';
when s1178 => state := s1179; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1179 => 			--14
	if (addfprdy = '1') then state := s1180;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1179; end if;
when s1180 => state := s1181; 	--15
	addfpsclr <= '0';
when s1181 => state := s1182; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1182 => 			--17
	if (addfprdy = '1') then state := s1183;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1182; end if;
when s1183 => state := s1184; 	--18
	addfpsclr <= '0';
when s1184 => state := s1185; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1185 => 			--20
	if (addfprdy = '1') then state := s1186;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1185; end if;
when s1186 => state := s1187; 	--21
	addfpsclr <= '0';
when s1187 => state := s1188; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (109, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1188 => state := s1189; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (156, 12)); -- offset LSB 108
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s1189 => state := s1190;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (157, 12)); -- offset MSB 109
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1190 => state := s1191; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1191 => 			--4
	if (fixed2floatrdy = '1') then state := s1192;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1191; end if;
when s1192 => state := s1193; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1193 => 			--6
	if (mulfprdy = '1') then state := s1194;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1193; end if;
when s1194 => state := s1195; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1195 => 			--8
	if (mulfprdy = '1') then state := s1196;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1195; end if;
when s1196 => state := s1197; 	--9
	mulfpsclr <= '0';
when s1197 => state := s1198; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1198 => 			--11
	if (mulfprdy = '1') then state := s1199;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1198; end if;
when s1199 => state := s1200; 	--12
	mulfpsclr <= '0';
when s1200 => state := s1201; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1201 => 			--14
	if (addfprdy = '1') then state := s1202;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1201; end if;
when s1202 => state := s1203; 	--15
	addfpsclr <= '0';
when s1203 => state := s1204; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1204 => 			--17
	if (addfprdy = '1') then state := s1205;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1204; end if;
when s1205 => state := s1206; 	--18
	addfpsclr <= '0';
when s1206 => state := s1207; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1207 => 			--20
	if (addfprdy = '1') then state := s1208;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1207; end if;
when s1208 => state := s1209; 	--21
	addfpsclr <= '0';
when s1209 => state := s1210; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (110, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1210 => state := s1211; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (158, 12)); -- offset LSB 110
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s1211 => state := s1212;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (159, 12)); -- offset MSB 111
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1212 => state := s1213; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1213 => 			--4
	if (fixed2floatrdy = '1') then state := s1214;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1213; end if;
when s1214 => state := s1215; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1215 => 			--6
	if (mulfprdy = '1') then state := s1216;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1215; end if;
when s1216 => state := s1217; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1217 => 			--8
	if (mulfprdy = '1') then state := s1218;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1217; end if;
when s1218 => state := s1219; 	--9
	mulfpsclr <= '0';
when s1219 => state := s1220; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1220 => 			--11
	if (mulfprdy = '1') then state := s1221;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1220; end if;
when s1221 => state := s1222; 	--12
	mulfpsclr <= '0';
when s1222 => state := s1223; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1223 => 			--14
	if (addfprdy = '1') then state := s1224;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1223; end if;
when s1224 => state := s1225; 	--15
	addfpsclr <= '0';
when s1225 => state := s1226; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1226 => 			--17
	if (addfprdy = '1') then state := s1227;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1226; end if;
when s1227 => state := s1228; 	--18
	addfpsclr <= '0';
when s1228 => state := s1229; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1229 => 			--20
	if (addfprdy = '1') then state := s1230;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1229; end if;
when s1230 => state := s1231; 	--21
	addfpsclr <= '0';
when s1231 => state := s1232; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (111, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1232 => state := s1233; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (160, 12)); -- offset LSB 112
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s1233 => state := s1234;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (161, 12)); -- offset MSB 113
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1234 => state := s1235; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1235 => 			--4
	if (fixed2floatrdy = '1') then state := s1236;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1235; end if;
when s1236 => state := s1237; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1237 => 			--6
	if (mulfprdy = '1') then state := s1238;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1237; end if;
when s1238 => state := s1239; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1239 => 			--8
	if (mulfprdy = '1') then state := s1240;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1239; end if;
when s1240 => state := s1241; 	--9
	mulfpsclr <= '0';
when s1241 => state := s1242; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1242 => 			--11
	if (mulfprdy = '1') then state := s1243;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1242; end if;
when s1243 => state := s1244; 	--12
	mulfpsclr <= '0';
when s1244 => state := s1245; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1245 => 			--14
	if (addfprdy = '1') then state := s1246;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1245; end if;
when s1246 => state := s1247; 	--15
	addfpsclr <= '0';
when s1247 => state := s1248; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1248 => 			--17
	if (addfprdy = '1') then state := s1249;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1248; end if;
when s1249 => state := s1250; 	--18
	addfpsclr <= '0';
when s1250 => state := s1251; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1251 => 			--20
	if (addfprdy = '1') then state := s1252;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1251; end if;
when s1252 => state := s1253; 	--21
	addfpsclr <= '0';
when s1253 => state := s1254; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (112, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1254 => state := s1255; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (162, 12)); -- offset LSB 114
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s1255 => state := s1256;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (163, 12)); -- offset MSB 115
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1256 => state := s1257; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1257 => 			--4
	if (fixed2floatrdy = '1') then state := s1258;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1257; end if;
when s1258 => state := s1259; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1259 => 			--6
	if (mulfprdy = '1') then state := s1260;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1259; end if;
when s1260 => state := s1261; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1261 => 			--8
	if (mulfprdy = '1') then state := s1262;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1261; end if;
when s1262 => state := s1263; 	--9
	mulfpsclr <= '0';
when s1263 => state := s1264; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1264 => 			--11
	if (mulfprdy = '1') then state := s1265;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1264; end if;
when s1265 => state := s1266; 	--12
	mulfpsclr <= '0';
when s1266 => state := s1267; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1267 => 			--14
	if (addfprdy = '1') then state := s1268;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1267; end if;
when s1268 => state := s1269; 	--15
	addfpsclr <= '0';
when s1269 => state := s1270; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1270 => 			--17
	if (addfprdy = '1') then state := s1271;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1270; end if;
when s1271 => state := s1272; 	--18
	addfpsclr <= '0';
when s1272 => state := s1273; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1273 => 			--20
	if (addfprdy = '1') then state := s1274;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1273; end if;
when s1274 => state := s1275; 	--21
	addfpsclr <= '0';
when s1275 => state := s1276; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (113, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1276 => state := s1277; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (164, 12)); -- offset LSB 116
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s1277 => state := s1278;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (165, 12)); -- offset MSB 117
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1278 => state := s1279; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1279 => 			--4
	if (fixed2floatrdy = '1') then state := s1280;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1279; end if;
when s1280 => state := s1281; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1281 => 			--6
	if (mulfprdy = '1') then state := s1282;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1281; end if;
when s1282 => state := s1283; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1283 => 			--8
	if (mulfprdy = '1') then state := s1284;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1283; end if;
when s1284 => state := s1285; 	--9
	mulfpsclr <= '0';
when s1285 => state := s1286; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1286 => 			--11
	if (mulfprdy = '1') then state := s1287;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1286; end if;
when s1287 => state := s1288; 	--12
	mulfpsclr <= '0';
when s1288 => state := s1289; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1289 => 			--14
	if (addfprdy = '1') then state := s1290;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1289; end if;
when s1290 => state := s1291; 	--15
	addfpsclr <= '0';
when s1291 => state := s1292; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1292 => 			--17
	if (addfprdy = '1') then state := s1293;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1292; end if;
when s1293 => state := s1294; 	--18
	addfpsclr <= '0';
when s1294 => state := s1295; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1295 => 			--20
	if (addfprdy = '1') then state := s1296;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1295; end if;
when s1296 => state := s1297; 	--21
	addfpsclr <= '0';
when s1297 => state := s1298; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (114, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1298 => state := s1299; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (166, 12)); -- offset LSB 118
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s1299 => state := s1300;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (167, 12)); -- offset MSB 119
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1300 => state := s1301; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1301 => 			--4
	if (fixed2floatrdy = '1') then state := s1302;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1301; end if;
when s1302 => state := s1303; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1303 => 			--6
	if (mulfprdy = '1') then state := s1304;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1303; end if;
when s1304 => state := s1305; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1305 => 			--8
	if (mulfprdy = '1') then state := s1306;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1305; end if;
when s1306 => state := s1307; 	--9
	mulfpsclr <= '0';
when s1307 => state := s1308; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1308 => 			--11
	if (mulfprdy = '1') then state := s1309;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1308; end if;
when s1309 => state := s1310; 	--12
	mulfpsclr <= '0';
when s1310 => state := s1311; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1311 => 			--14
	if (addfprdy = '1') then state := s1312;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1311; end if;
when s1312 => state := s1313; 	--15
	addfpsclr <= '0';
when s1313 => state := s1314; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1314 => 			--17
	if (addfprdy = '1') then state := s1315;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1314; end if;
when s1315 => state := s1316; 	--18
	addfpsclr <= '0';
when s1316 => state := s1317; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1317 => 			--20
	if (addfprdy = '1') then state := s1318;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1317; end if;
when s1318 => state := s1319; 	--21
	addfpsclr <= '0';
when s1319 => state := s1320; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (115, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1320 => state := s1321; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (168, 12)); -- offset LSB 120
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s1321 => state := s1322;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (169, 12)); -- offset MSB 121
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1322 => state := s1323; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1323 => 			--4
	if (fixed2floatrdy = '1') then state := s1324;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1323; end if;
when s1324 => state := s1325; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1325 => 			--6
	if (mulfprdy = '1') then state := s1326;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1325; end if;
when s1326 => state := s1327; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1327 => 			--8
	if (mulfprdy = '1') then state := s1328;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1327; end if;
when s1328 => state := s1329; 	--9
	mulfpsclr <= '0';
when s1329 => state := s1330; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1330 => 			--11
	if (mulfprdy = '1') then state := s1331;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1330; end if;
when s1331 => state := s1332; 	--12
	mulfpsclr <= '0';
when s1332 => state := s1333; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1333 => 			--14
	if (addfprdy = '1') then state := s1334;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1333; end if;
when s1334 => state := s1335; 	--15
	addfpsclr <= '0';
when s1335 => state := s1336; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1336 => 			--17
	if (addfprdy = '1') then state := s1337;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1336; end if;
when s1337 => state := s1338; 	--18
	addfpsclr <= '0';
when s1338 => state := s1339; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1339 => 			--20
	if (addfprdy = '1') then state := s1340;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1339; end if;
when s1340 => state := s1341; 	--21
	addfpsclr <= '0';
when s1341 => state := s1342; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (116, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1342 => state := s1343; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (170, 12)); -- offset LSB 122
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s1343 => state := s1344;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (171, 12)); -- offset MSB 123
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1344 => state := s1345; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1345 => 			--4
	if (fixed2floatrdy = '1') then state := s1346;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1345; end if;
when s1346 => state := s1347; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1347 => 			--6
	if (mulfprdy = '1') then state := s1348;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1347; end if;
when s1348 => state := s1349; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1349 => 			--8
	if (mulfprdy = '1') then state := s1350;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1349; end if;
when s1350 => state := s1351; 	--9
	mulfpsclr <= '0';
when s1351 => state := s1352; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1352 => 			--11
	if (mulfprdy = '1') then state := s1353;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1352; end if;
when s1353 => state := s1354; 	--12
	mulfpsclr <= '0';
when s1354 => state := s1355; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1355 => 			--14
	if (addfprdy = '1') then state := s1356;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1355; end if;
when s1356 => state := s1357; 	--15
	addfpsclr <= '0';
when s1357 => state := s1358; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1358 => 			--17
	if (addfprdy = '1') then state := s1359;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1358; end if;
when s1359 => state := s1360; 	--18
	addfpsclr <= '0';
when s1360 => state := s1361; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1361 => 			--20
	if (addfprdy = '1') then state := s1362;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1361; end if;
when s1362 => state := s1363; 	--21
	addfpsclr <= '0';
when s1363 => state := s1364; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (117, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1364 => state := s1365; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (172, 12)); -- offset LSB 124
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s1365 => state := s1366;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (173, 12)); -- offset MSB 125
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1366 => state := s1367; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1367 => 			--4
	if (fixed2floatrdy = '1') then state := s1368;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1367; end if;
when s1368 => state := s1369; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1369 => 			--6
	if (mulfprdy = '1') then state := s1370;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1369; end if;
when s1370 => state := s1371; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1371 => 			--8
	if (mulfprdy = '1') then state := s1372;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1371; end if;
when s1372 => state := s1373; 	--9
	mulfpsclr <= '0';
when s1373 => state := s1374; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1374 => 			--11
	if (mulfprdy = '1') then state := s1375;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1374; end if;
when s1375 => state := s1376; 	--12
	mulfpsclr <= '0';
when s1376 => state := s1377; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1377 => 			--14
	if (addfprdy = '1') then state := s1378;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1377; end if;
when s1378 => state := s1379; 	--15
	addfpsclr <= '0';
when s1379 => state := s1380; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1380 => 			--17
	if (addfprdy = '1') then state := s1381;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1380; end if;
when s1381 => state := s1382; 	--18
	addfpsclr <= '0';
when s1382 => state := s1383; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1383 => 			--20
	if (addfprdy = '1') then state := s1384;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1383; end if;
when s1384 => state := s1385; 	--21
	addfpsclr <= '0';
when s1385 => state := s1386; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (118, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1386 => state := s1387; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (174, 12)); -- offset LSB 126
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s1387 => state := s1388;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (175, 12)); -- offset MSB 127
	addra <= std_logic_vector (to_unsigned (1, 10)); -- OCCrowI 1
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1388 => state := s1389; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1389 => 			--4
	if (fixed2floatrdy = '1') then state := s1390;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1389; end if;
when s1390 => state := s1391; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1391 => 			--6
	if (mulfprdy = '1') then state := s1392;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1391; end if;
when s1392 => state := s1393; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1393 => 			--8
	if (mulfprdy = '1') then state := s1394;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1393; end if;
when s1394 => state := s1395; 	--9
	mulfpsclr <= '0';
when s1395 => state := s1396; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1396 => 			--11
	if (mulfprdy = '1') then state := s1397;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1396; end if;
when s1397 => state := s1398; 	--12
	mulfpsclr <= '0';
when s1398 => state := s1399; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1399 => 			--14
	if (addfprdy = '1') then state := s1400;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1399; end if;
when s1400 => state := s1401; 	--15
	addfpsclr <= '0';
when s1401 => state := s1402; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1402 => 			--17
	if (addfprdy = '1') then state := s1403;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1402; end if;
when s1403 => state := s1404; 	--18
	addfpsclr <= '0';
when s1404 => state := s1405; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1405 => 			--20
	if (addfprdy = '1') then state := s1406;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1405; end if;
when s1406 => state := s1407; 	--21
	addfpsclr <= '0';
when s1407 => state := s1408; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (119, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1408 => state := s1409; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (176, 12)); -- offset LSB 128
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s1409 => state := s1410;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (177, 12)); -- offset MSB 129
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1410 => state := s1411; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1411 => 			--4
	if (fixed2floatrdy = '1') then state := s1412;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1411; end if;
when s1412 => state := s1413; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1413 => 			--6
	if (mulfprdy = '1') then state := s1414;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1413; end if;
when s1414 => state := s1415; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1415 => 			--8
	if (mulfprdy = '1') then state := s1416;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1415; end if;
when s1416 => state := s1417; 	--9
	mulfpsclr <= '0';
when s1417 => state := s1418; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1418 => 			--11
	if (mulfprdy = '1') then state := s1419;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1418; end if;
when s1419 => state := s1420; 	--12
	mulfpsclr <= '0';
when s1420 => state := s1421; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1421 => 			--14
	if (addfprdy = '1') then state := s1422;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1421; end if;
when s1422 => state := s1423; 	--15
	addfpsclr <= '0';
when s1423 => state := s1424; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1424 => 			--17
	if (addfprdy = '1') then state := s1425;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1424; end if;
when s1425 => state := s1426; 	--18
	addfpsclr <= '0';
when s1426 => state := s1427; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1427 => 			--20
	if (addfprdy = '1') then state := s1428;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1427; end if;
when s1428 => state := s1429; 	--21
	addfpsclr <= '0';
when s1429 => state := s1430; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (120, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1430 => state := s1431; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (178, 12)); -- offset LSB 130
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s1431 => state := s1432;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (179, 12)); -- offset MSB 131
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1432 => state := s1433; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1433 => 			--4
	if (fixed2floatrdy = '1') then state := s1434;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1433; end if;
when s1434 => state := s1435; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1435 => 			--6
	if (mulfprdy = '1') then state := s1436;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1435; end if;
when s1436 => state := s1437; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1437 => 			--8
	if (mulfprdy = '1') then state := s1438;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1437; end if;
when s1438 => state := s1439; 	--9
	mulfpsclr <= '0';
when s1439 => state := s1440; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1440 => 			--11
	if (mulfprdy = '1') then state := s1441;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1440; end if;
when s1441 => state := s1442; 	--12
	mulfpsclr <= '0';
when s1442 => state := s1443; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1443 => 			--14
	if (addfprdy = '1') then state := s1444;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1443; end if;
when s1444 => state := s1445; 	--15
	addfpsclr <= '0';
when s1445 => state := s1446; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1446 => 			--17
	if (addfprdy = '1') then state := s1447;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1446; end if;
when s1447 => state := s1448; 	--18
	addfpsclr <= '0';
when s1448 => state := s1449; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1449 => 			--20
	if (addfprdy = '1') then state := s1450;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1449; end if;
when s1450 => state := s1451; 	--21
	addfpsclr <= '0';
when s1451 => state := s1452; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (121, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1452 => state := s1453; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (180, 12)); -- offset LSB 132
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s1453 => state := s1454;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (181, 12)); -- offset MSB 133
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1454 => state := s1455; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1455 => 			--4
	if (fixed2floatrdy = '1') then state := s1456;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1455; end if;
when s1456 => state := s1457; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1457 => 			--6
	if (mulfprdy = '1') then state := s1458;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1457; end if;
when s1458 => state := s1459; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1459 => 			--8
	if (mulfprdy = '1') then state := s1460;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1459; end if;
when s1460 => state := s1461; 	--9
	mulfpsclr <= '0';
when s1461 => state := s1462; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1462 => 			--11
	if (mulfprdy = '1') then state := s1463;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1462; end if;
when s1463 => state := s1464; 	--12
	mulfpsclr <= '0';
when s1464 => state := s1465; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1465 => 			--14
	if (addfprdy = '1') then state := s1466;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1465; end if;
when s1466 => state := s1467; 	--15
	addfpsclr <= '0';
when s1467 => state := s1468; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1468 => 			--17
	if (addfprdy = '1') then state := s1469;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1468; end if;
when s1469 => state := s1470; 	--18
	addfpsclr <= '0';
when s1470 => state := s1471; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1471 => 			--20
	if (addfprdy = '1') then state := s1472;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1471; end if;
when s1472 => state := s1473; 	--21
	addfpsclr <= '0';
when s1473 => state := s1474; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (122, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1474 => state := s1475; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (182, 12)); -- offset LSB 134
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s1475 => state := s1476;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (183, 12)); -- offset MSB 135
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1476 => state := s1477; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1477 => 			--4
	if (fixed2floatrdy = '1') then state := s1478;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1477; end if;
when s1478 => state := s1479; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1479 => 			--6
	if (mulfprdy = '1') then state := s1480;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1479; end if;
when s1480 => state := s1481; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1481 => 			--8
	if (mulfprdy = '1') then state := s1482;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1481; end if;
when s1482 => state := s1483; 	--9
	mulfpsclr <= '0';
when s1483 => state := s1484; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1484 => 			--11
	if (mulfprdy = '1') then state := s1485;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1484; end if;
when s1485 => state := s1486; 	--12
	mulfpsclr <= '0';
when s1486 => state := s1487; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1487 => 			--14
	if (addfprdy = '1') then state := s1488;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1487; end if;
when s1488 => state := s1489; 	--15
	addfpsclr <= '0';
when s1489 => state := s1490; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1490 => 			--17
	if (addfprdy = '1') then state := s1491;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1490; end if;
when s1491 => state := s1492; 	--18
	addfpsclr <= '0';
when s1492 => state := s1493; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1493 => 			--20
	if (addfprdy = '1') then state := s1494;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1493; end if;
when s1494 => state := s1495; 	--21
	addfpsclr <= '0';
when s1495 => state := s1496; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (123, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1496 => state := s1497; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (184, 12)); -- offset LSB 136
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s1497 => state := s1498;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (185, 12)); -- offset MSB 137
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1498 => state := s1499; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1499 => 			--4
	if (fixed2floatrdy = '1') then state := s1500;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1499; end if;
when s1500 => state := s1501; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1501 => 			--6
	if (mulfprdy = '1') then state := s1502;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1501; end if;
when s1502 => state := s1503; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1503 => 			--8
	if (mulfprdy = '1') then state := s1504;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1503; end if;
when s1504 => state := s1505; 	--9
	mulfpsclr <= '0';
when s1505 => state := s1506; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1506 => 			--11
	if (mulfprdy = '1') then state := s1507;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1506; end if;
when s1507 => state := s1508; 	--12
	mulfpsclr <= '0';
when s1508 => state := s1509; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1509 => 			--14
	if (addfprdy = '1') then state := s1510;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1509; end if;
when s1510 => state := s1511; 	--15
	addfpsclr <= '0';
when s1511 => state := s1512; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1512 => 			--17
	if (addfprdy = '1') then state := s1513;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1512; end if;
when s1513 => state := s1514; 	--18
	addfpsclr <= '0';
when s1514 => state := s1515; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1515 => 			--20
	if (addfprdy = '1') then state := s1516;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1515; end if;
when s1516 => state := s1517; 	--21
	addfpsclr <= '0';
when s1517 => state := s1518; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (124, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1518 => state := s1519; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (186, 12)); -- offset LSB 138
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s1519 => state := s1520;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (187, 12)); -- offset MSB 139
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1520 => state := s1521; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1521 => 			--4
	if (fixed2floatrdy = '1') then state := s1522;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1521; end if;
when s1522 => state := s1523; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1523 => 			--6
	if (mulfprdy = '1') then state := s1524;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1523; end if;
when s1524 => state := s1525; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1525 => 			--8
	if (mulfprdy = '1') then state := s1526;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1525; end if;
when s1526 => state := s1527; 	--9
	mulfpsclr <= '0';
when s1527 => state := s1528; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1528 => 			--11
	if (mulfprdy = '1') then state := s1529;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1528; end if;
when s1529 => state := s1530; 	--12
	mulfpsclr <= '0';
when s1530 => state := s1531; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1531 => 			--14
	if (addfprdy = '1') then state := s1532;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1531; end if;
when s1532 => state := s1533; 	--15
	addfpsclr <= '0';
when s1533 => state := s1534; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1534 => 			--17
	if (addfprdy = '1') then state := s1535;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1534; end if;
when s1535 => state := s1536; 	--18
	addfpsclr <= '0';
when s1536 => state := s1537; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1537 => 			--20
	if (addfprdy = '1') then state := s1538;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1537; end if;
when s1538 => state := s1539; 	--21
	addfpsclr <= '0';
when s1539 => state := s1540; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (125, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1540 => state := s1541; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (188, 12)); -- offset LSB 140
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s1541 => state := s1542;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (189, 12)); -- offset MSB 141
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1542 => state := s1543; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1543 => 			--4
	if (fixed2floatrdy = '1') then state := s1544;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1543; end if;
when s1544 => state := s1545; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1545 => 			--6
	if (mulfprdy = '1') then state := s1546;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1545; end if;
when s1546 => state := s1547; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1547 => 			--8
	if (mulfprdy = '1') then state := s1548;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1547; end if;
when s1548 => state := s1549; 	--9
	mulfpsclr <= '0';
when s1549 => state := s1550; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1550 => 			--11
	if (mulfprdy = '1') then state := s1551;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1550; end if;
when s1551 => state := s1552; 	--12
	mulfpsclr <= '0';
when s1552 => state := s1553; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1553 => 			--14
	if (addfprdy = '1') then state := s1554;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1553; end if;
when s1554 => state := s1555; 	--15
	addfpsclr <= '0';
when s1555 => state := s1556; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1556 => 			--17
	if (addfprdy = '1') then state := s1557;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1556; end if;
when s1557 => state := s1558; 	--18
	addfpsclr <= '0';
when s1558 => state := s1559; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1559 => 			--20
	if (addfprdy = '1') then state := s1560;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1559; end if;
when s1560 => state := s1561; 	--21
	addfpsclr <= '0';
when s1561 => state := s1562; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (126, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1562 => state := s1563; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (190, 12)); -- offset LSB 142
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s1563 => state := s1564;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (191, 12)); -- offset MSB 143
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1564 => state := s1565; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1565 => 			--4
	if (fixed2floatrdy = '1') then state := s1566;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1565; end if;
when s1566 => state := s1567; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1567 => 			--6
	if (mulfprdy = '1') then state := s1568;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1567; end if;
when s1568 => state := s1569; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1569 => 			--8
	if (mulfprdy = '1') then state := s1570;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1569; end if;
when s1570 => state := s1571; 	--9
	mulfpsclr <= '0';
when s1571 => state := s1572; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1572 => 			--11
	if (mulfprdy = '1') then state := s1573;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1572; end if;
when s1573 => state := s1574; 	--12
	mulfpsclr <= '0';
when s1574 => state := s1575; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1575 => 			--14
	if (addfprdy = '1') then state := s1576;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1575; end if;
when s1576 => state := s1577; 	--15
	addfpsclr <= '0';
when s1577 => state := s1578; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1578 => 			--17
	if (addfprdy = '1') then state := s1579;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1578; end if;
when s1579 => state := s1580; 	--18
	addfpsclr <= '0';
when s1580 => state := s1581; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1581 => 			--20
	if (addfprdy = '1') then state := s1582;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1581; end if;
when s1582 => state := s1583; 	--21
	addfpsclr <= '0';
when s1583 => state := s1584; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (127, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1584 => state := s1585; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (192, 12)); -- offset LSB 144
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s1585 => state := s1586;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (193, 12)); -- offset MSB 145
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1586 => state := s1587; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1587 => 			--4
	if (fixed2floatrdy = '1') then state := s1588;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1587; end if;
when s1588 => state := s1589; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1589 => 			--6
	if (mulfprdy = '1') then state := s1590;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1589; end if;
when s1590 => state := s1591; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1591 => 			--8
	if (mulfprdy = '1') then state := s1592;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1591; end if;
when s1592 => state := s1593; 	--9
	mulfpsclr <= '0';
when s1593 => state := s1594; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1594 => 			--11
	if (mulfprdy = '1') then state := s1595;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1594; end if;
when s1595 => state := s1596; 	--12
	mulfpsclr <= '0';
when s1596 => state := s1597; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1597 => 			--14
	if (addfprdy = '1') then state := s1598;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1597; end if;
when s1598 => state := s1599; 	--15
	addfpsclr <= '0';
when s1599 => state := s1600; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1600 => 			--17
	if (addfprdy = '1') then state := s1601;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1600; end if;
when s1601 => state := s1602; 	--18
	addfpsclr <= '0';
when s1602 => state := s1603; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1603 => 			--20
	if (addfprdy = '1') then state := s1604;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1603; end if;
when s1604 => state := s1605; 	--21
	addfpsclr <= '0';
when s1605 => state := s1606; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (128, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1606 => state := s1607; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (194, 12)); -- offset LSB 146
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s1607 => state := s1608;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (195, 12)); -- offset MSB 147
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1608 => state := s1609; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1609 => 			--4
	if (fixed2floatrdy = '1') then state := s1610;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1609; end if;
when s1610 => state := s1611; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1611 => 			--6
	if (mulfprdy = '1') then state := s1612;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1611; end if;
when s1612 => state := s1613; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1613 => 			--8
	if (mulfprdy = '1') then state := s1614;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1613; end if;
when s1614 => state := s1615; 	--9
	mulfpsclr <= '0';
when s1615 => state := s1616; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1616 => 			--11
	if (mulfprdy = '1') then state := s1617;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1616; end if;
when s1617 => state := s1618; 	--12
	mulfpsclr <= '0';
when s1618 => state := s1619; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1619 => 			--14
	if (addfprdy = '1') then state := s1620;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1619; end if;
when s1620 => state := s1621; 	--15
	addfpsclr <= '0';
when s1621 => state := s1622; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1622 => 			--17
	if (addfprdy = '1') then state := s1623;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1622; end if;
when s1623 => state := s1624; 	--18
	addfpsclr <= '0';
when s1624 => state := s1625; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1625 => 			--20
	if (addfprdy = '1') then state := s1626;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1625; end if;
when s1626 => state := s1627; 	--21
	addfpsclr <= '0';
when s1627 => state := s1628; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (129, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1628 => state := s1629; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (196, 12)); -- offset LSB 148
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s1629 => state := s1630;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (197, 12)); -- offset MSB 149
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1630 => state := s1631; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1631 => 			--4
	if (fixed2floatrdy = '1') then state := s1632;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1631; end if;
when s1632 => state := s1633; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1633 => 			--6
	if (mulfprdy = '1') then state := s1634;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1633; end if;
when s1634 => state := s1635; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1635 => 			--8
	if (mulfprdy = '1') then state := s1636;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1635; end if;
when s1636 => state := s1637; 	--9
	mulfpsclr <= '0';
when s1637 => state := s1638; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1638 => 			--11
	if (mulfprdy = '1') then state := s1639;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1638; end if;
when s1639 => state := s1640; 	--12
	mulfpsclr <= '0';
when s1640 => state := s1641; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1641 => 			--14
	if (addfprdy = '1') then state := s1642;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1641; end if;
when s1642 => state := s1643; 	--15
	addfpsclr <= '0';
when s1643 => state := s1644; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1644 => 			--17
	if (addfprdy = '1') then state := s1645;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1644; end if;
when s1645 => state := s1646; 	--18
	addfpsclr <= '0';
when s1646 => state := s1647; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1647 => 			--20
	if (addfprdy = '1') then state := s1648;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1647; end if;
when s1648 => state := s1649; 	--21
	addfpsclr <= '0';
when s1649 => state := s1650; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (130, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1650 => state := s1651; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (198, 12)); -- offset LSB 150
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s1651 => state := s1652;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (199, 12)); -- offset MSB 151
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1652 => state := s1653; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1653 => 			--4
	if (fixed2floatrdy = '1') then state := s1654;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1653; end if;
when s1654 => state := s1655; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1655 => 			--6
	if (mulfprdy = '1') then state := s1656;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1655; end if;
when s1656 => state := s1657; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1657 => 			--8
	if (mulfprdy = '1') then state := s1658;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1657; end if;
when s1658 => state := s1659; 	--9
	mulfpsclr <= '0';
when s1659 => state := s1660; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1660 => 			--11
	if (mulfprdy = '1') then state := s1661;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1660; end if;
when s1661 => state := s1662; 	--12
	mulfpsclr <= '0';
when s1662 => state := s1663; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1663 => 			--14
	if (addfprdy = '1') then state := s1664;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1663; end if;
when s1664 => state := s1665; 	--15
	addfpsclr <= '0';
when s1665 => state := s1666; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1666 => 			--17
	if (addfprdy = '1') then state := s1667;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1666; end if;
when s1667 => state := s1668; 	--18
	addfpsclr <= '0';
when s1668 => state := s1669; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1669 => 			--20
	if (addfprdy = '1') then state := s1670;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1669; end if;
when s1670 => state := s1671; 	--21
	addfpsclr <= '0';
when s1671 => state := s1672; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (131, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1672 => state := s1673; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (200, 12)); -- offset LSB 152
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s1673 => state := s1674;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (201, 12)); -- offset MSB 153
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1674 => state := s1675; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1675 => 			--4
	if (fixed2floatrdy = '1') then state := s1676;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1675; end if;
when s1676 => state := s1677; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1677 => 			--6
	if (mulfprdy = '1') then state := s1678;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1677; end if;
when s1678 => state := s1679; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1679 => 			--8
	if (mulfprdy = '1') then state := s1680;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1679; end if;
when s1680 => state := s1681; 	--9
	mulfpsclr <= '0';
when s1681 => state := s1682; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1682 => 			--11
	if (mulfprdy = '1') then state := s1683;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1682; end if;
when s1683 => state := s1684; 	--12
	mulfpsclr <= '0';
when s1684 => state := s1685; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1685 => 			--14
	if (addfprdy = '1') then state := s1686;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1685; end if;
when s1686 => state := s1687; 	--15
	addfpsclr <= '0';
when s1687 => state := s1688; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1688 => 			--17
	if (addfprdy = '1') then state := s1689;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1688; end if;
when s1689 => state := s1690; 	--18
	addfpsclr <= '0';
when s1690 => state := s1691; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1691 => 			--20
	if (addfprdy = '1') then state := s1692;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1691; end if;
when s1692 => state := s1693; 	--21
	addfpsclr <= '0';
when s1693 => state := s1694; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (132, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1694 => state := s1695; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (202, 12)); -- offset LSB 154
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s1695 => state := s1696;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (203, 12)); -- offset MSB 155
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1696 => state := s1697; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1697 => 			--4
	if (fixed2floatrdy = '1') then state := s1698;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1697; end if;
when s1698 => state := s1699; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1699 => 			--6
	if (mulfprdy = '1') then state := s1700;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1699; end if;
when s1700 => state := s1701; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1701 => 			--8
	if (mulfprdy = '1') then state := s1702;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1701; end if;
when s1702 => state := s1703; 	--9
	mulfpsclr <= '0';
when s1703 => state := s1704; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1704 => 			--11
	if (mulfprdy = '1') then state := s1705;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1704; end if;
when s1705 => state := s1706; 	--12
	mulfpsclr <= '0';
when s1706 => state := s1707; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1707 => 			--14
	if (addfprdy = '1') then state := s1708;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1707; end if;
when s1708 => state := s1709; 	--15
	addfpsclr <= '0';
when s1709 => state := s1710; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1710 => 			--17
	if (addfprdy = '1') then state := s1711;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1710; end if;
when s1711 => state := s1712; 	--18
	addfpsclr <= '0';
when s1712 => state := s1713; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1713 => 			--20
	if (addfprdy = '1') then state := s1714;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1713; end if;
when s1714 => state := s1715; 	--21
	addfpsclr <= '0';
when s1715 => state := s1716; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (133, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1716 => state := s1717; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (204, 12)); -- offset LSB 156
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s1717 => state := s1718;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (205, 12)); -- offset MSB 157
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1718 => state := s1719; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1719 => 			--4
	if (fixed2floatrdy = '1') then state := s1720;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1719; end if;
when s1720 => state := s1721; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1721 => 			--6
	if (mulfprdy = '1') then state := s1722;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1721; end if;
when s1722 => state := s1723; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1723 => 			--8
	if (mulfprdy = '1') then state := s1724;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1723; end if;
when s1724 => state := s1725; 	--9
	mulfpsclr <= '0';
when s1725 => state := s1726; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1726 => 			--11
	if (mulfprdy = '1') then state := s1727;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1726; end if;
when s1727 => state := s1728; 	--12
	mulfpsclr <= '0';
when s1728 => state := s1729; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1729 => 			--14
	if (addfprdy = '1') then state := s1730;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1729; end if;
when s1730 => state := s1731; 	--15
	addfpsclr <= '0';
when s1731 => state := s1732; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1732 => 			--17
	if (addfprdy = '1') then state := s1733;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1732; end if;
when s1733 => state := s1734; 	--18
	addfpsclr <= '0';
when s1734 => state := s1735; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1735 => 			--20
	if (addfprdy = '1') then state := s1736;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1735; end if;
when s1736 => state := s1737; 	--21
	addfpsclr <= '0';
when s1737 => state := s1738; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (134, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1738 => state := s1739; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (206, 12)); -- offset LSB 158
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s1739 => state := s1740;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (207, 12)); -- offset MSB 159
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1740 => state := s1741; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1741 => 			--4
	if (fixed2floatrdy = '1') then state := s1742;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1741; end if;
when s1742 => state := s1743; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1743 => 			--6
	if (mulfprdy = '1') then state := s1744;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1743; end if;
when s1744 => state := s1745; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1745 => 			--8
	if (mulfprdy = '1') then state := s1746;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1745; end if;
when s1746 => state := s1747; 	--9
	mulfpsclr <= '0';
when s1747 => state := s1748; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1748 => 			--11
	if (mulfprdy = '1') then state := s1749;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1748; end if;
when s1749 => state := s1750; 	--12
	mulfpsclr <= '0';
when s1750 => state := s1751; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1751 => 			--14
	if (addfprdy = '1') then state := s1752;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1751; end if;
when s1752 => state := s1753; 	--15
	addfpsclr <= '0';
when s1753 => state := s1754; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1754 => 			--17
	if (addfprdy = '1') then state := s1755;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1754; end if;
when s1755 => state := s1756; 	--18
	addfpsclr <= '0';
when s1756 => state := s1757; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1757 => 			--20
	if (addfprdy = '1') then state := s1758;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1757; end if;
when s1758 => state := s1759; 	--21
	addfpsclr <= '0';
when s1759 => state := s1760; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (135, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1760 => state := s1761; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (208, 12)); -- offset LSB 160
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s1761 => state := s1762;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (209, 12)); -- offset MSB 161
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1762 => state := s1763; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1763 => 			--4
	if (fixed2floatrdy = '1') then state := s1764;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1763; end if;
when s1764 => state := s1765; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1765 => 			--6
	if (mulfprdy = '1') then state := s1766;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1765; end if;
when s1766 => state := s1767; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1767 => 			--8
	if (mulfprdy = '1') then state := s1768;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1767; end if;
when s1768 => state := s1769; 	--9
	mulfpsclr <= '0';
when s1769 => state := s1770; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1770 => 			--11
	if (mulfprdy = '1') then state := s1771;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1770; end if;
when s1771 => state := s1772; 	--12
	mulfpsclr <= '0';
when s1772 => state := s1773; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1773 => 			--14
	if (addfprdy = '1') then state := s1774;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1773; end if;
when s1774 => state := s1775; 	--15
	addfpsclr <= '0';
when s1775 => state := s1776; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1776 => 			--17
	if (addfprdy = '1') then state := s1777;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1776; end if;
when s1777 => state := s1778; 	--18
	addfpsclr <= '0';
when s1778 => state := s1779; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1779 => 			--20
	if (addfprdy = '1') then state := s1780;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1779; end if;
when s1780 => state := s1781; 	--21
	addfpsclr <= '0';
when s1781 => state := s1782; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (136, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1782 => state := s1783; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (210, 12)); -- offset LSB 162
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s1783 => state := s1784;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (211, 12)); -- offset MSB 163
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1784 => state := s1785; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1785 => 			--4
	if (fixed2floatrdy = '1') then state := s1786;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1785; end if;
when s1786 => state := s1787; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1787 => 			--6
	if (mulfprdy = '1') then state := s1788;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1787; end if;
when s1788 => state := s1789; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1789 => 			--8
	if (mulfprdy = '1') then state := s1790;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1789; end if;
when s1790 => state := s1791; 	--9
	mulfpsclr <= '0';
when s1791 => state := s1792; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1792 => 			--11
	if (mulfprdy = '1') then state := s1793;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1792; end if;
when s1793 => state := s1794; 	--12
	mulfpsclr <= '0';
when s1794 => state := s1795; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1795 => 			--14
	if (addfprdy = '1') then state := s1796;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1795; end if;
when s1796 => state := s1797; 	--15
	addfpsclr <= '0';
when s1797 => state := s1798; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1798 => 			--17
	if (addfprdy = '1') then state := s1799;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1798; end if;
when s1799 => state := s1800; 	--18
	addfpsclr <= '0';
when s1800 => state := s1801; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1801 => 			--20
	if (addfprdy = '1') then state := s1802;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1801; end if;
when s1802 => state := s1803; 	--21
	addfpsclr <= '0';
when s1803 => state := s1804; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (137, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1804 => state := s1805; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (212, 12)); -- offset LSB 164
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s1805 => state := s1806;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (213, 12)); -- offset MSB 165
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1806 => state := s1807; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1807 => 			--4
	if (fixed2floatrdy = '1') then state := s1808;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1807; end if;
when s1808 => state := s1809; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1809 => 			--6
	if (mulfprdy = '1') then state := s1810;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1809; end if;
when s1810 => state := s1811; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1811 => 			--8
	if (mulfprdy = '1') then state := s1812;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1811; end if;
when s1812 => state := s1813; 	--9
	mulfpsclr <= '0';
when s1813 => state := s1814; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1814 => 			--11
	if (mulfprdy = '1') then state := s1815;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1814; end if;
when s1815 => state := s1816; 	--12
	mulfpsclr <= '0';
when s1816 => state := s1817; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1817 => 			--14
	if (addfprdy = '1') then state := s1818;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1817; end if;
when s1818 => state := s1819; 	--15
	addfpsclr <= '0';
when s1819 => state := s1820; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1820 => 			--17
	if (addfprdy = '1') then state := s1821;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1820; end if;
when s1821 => state := s1822; 	--18
	addfpsclr <= '0';
when s1822 => state := s1823; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1823 => 			--20
	if (addfprdy = '1') then state := s1824;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1823; end if;
when s1824 => state := s1825; 	--21
	addfpsclr <= '0';
when s1825 => state := s1826; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (138, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1826 => state := s1827; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (214, 12)); -- offset LSB 166
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s1827 => state := s1828;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (215, 12)); -- offset MSB 167
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1828 => state := s1829; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1829 => 			--4
	if (fixed2floatrdy = '1') then state := s1830;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1829; end if;
when s1830 => state := s1831; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1831 => 			--6
	if (mulfprdy = '1') then state := s1832;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1831; end if;
when s1832 => state := s1833; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1833 => 			--8
	if (mulfprdy = '1') then state := s1834;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1833; end if;
when s1834 => state := s1835; 	--9
	mulfpsclr <= '0';
when s1835 => state := s1836; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1836 => 			--11
	if (mulfprdy = '1') then state := s1837;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1836; end if;
when s1837 => state := s1838; 	--12
	mulfpsclr <= '0';
when s1838 => state := s1839; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1839 => 			--14
	if (addfprdy = '1') then state := s1840;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1839; end if;
when s1840 => state := s1841; 	--15
	addfpsclr <= '0';
when s1841 => state := s1842; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1842 => 			--17
	if (addfprdy = '1') then state := s1843;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1842; end if;
when s1843 => state := s1844; 	--18
	addfpsclr <= '0';
when s1844 => state := s1845; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1845 => 			--20
	if (addfprdy = '1') then state := s1846;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1845; end if;
when s1846 => state := s1847; 	--21
	addfpsclr <= '0';
when s1847 => state := s1848; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (139, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1848 => state := s1849; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (216, 12)); -- offset LSB 168
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s1849 => state := s1850;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (217, 12)); -- offset MSB 169
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1850 => state := s1851; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1851 => 			--4
	if (fixed2floatrdy = '1') then state := s1852;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1851; end if;
when s1852 => state := s1853; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1853 => 			--6
	if (mulfprdy = '1') then state := s1854;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1853; end if;
when s1854 => state := s1855; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1855 => 			--8
	if (mulfprdy = '1') then state := s1856;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1855; end if;
when s1856 => state := s1857; 	--9
	mulfpsclr <= '0';
when s1857 => state := s1858; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1858 => 			--11
	if (mulfprdy = '1') then state := s1859;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1858; end if;
when s1859 => state := s1860; 	--12
	mulfpsclr <= '0';
when s1860 => state := s1861; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1861 => 			--14
	if (addfprdy = '1') then state := s1862;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1861; end if;
when s1862 => state := s1863; 	--15
	addfpsclr <= '0';
when s1863 => state := s1864; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1864 => 			--17
	if (addfprdy = '1') then state := s1865;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1864; end if;
when s1865 => state := s1866; 	--18
	addfpsclr <= '0';
when s1866 => state := s1867; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1867 => 			--20
	if (addfprdy = '1') then state := s1868;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1867; end if;
when s1868 => state := s1869; 	--21
	addfpsclr <= '0';
when s1869 => state := s1870; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (140, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1870 => state := s1871; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (218, 12)); -- offset LSB 170
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s1871 => state := s1872;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (219, 12)); -- offset MSB 171
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1872 => state := s1873; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1873 => 			--4
	if (fixed2floatrdy = '1') then state := s1874;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1873; end if;
when s1874 => state := s1875; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1875 => 			--6
	if (mulfprdy = '1') then state := s1876;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1875; end if;
when s1876 => state := s1877; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1877 => 			--8
	if (mulfprdy = '1') then state := s1878;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1877; end if;
when s1878 => state := s1879; 	--9
	mulfpsclr <= '0';
when s1879 => state := s1880; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1880 => 			--11
	if (mulfprdy = '1') then state := s1881;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1880; end if;
when s1881 => state := s1882; 	--12
	mulfpsclr <= '0';
when s1882 => state := s1883; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1883 => 			--14
	if (addfprdy = '1') then state := s1884;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1883; end if;
when s1884 => state := s1885; 	--15
	addfpsclr <= '0';
when s1885 => state := s1886; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1886 => 			--17
	if (addfprdy = '1') then state := s1887;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1886; end if;
when s1887 => state := s1888; 	--18
	addfpsclr <= '0';
when s1888 => state := s1889; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1889 => 			--20
	if (addfprdy = '1') then state := s1890;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1889; end if;
when s1890 => state := s1891; 	--21
	addfpsclr <= '0';
when s1891 => state := s1892; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (141, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1892 => state := s1893; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (220, 12)); -- offset LSB 172
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s1893 => state := s1894;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (221, 12)); -- offset MSB 173
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1894 => state := s1895; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1895 => 			--4
	if (fixed2floatrdy = '1') then state := s1896;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1895; end if;
when s1896 => state := s1897; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1897 => 			--6
	if (mulfprdy = '1') then state := s1898;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1897; end if;
when s1898 => state := s1899; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1899 => 			--8
	if (mulfprdy = '1') then state := s1900;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1899; end if;
when s1900 => state := s1901; 	--9
	mulfpsclr <= '0';
when s1901 => state := s1902; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1902 => 			--11
	if (mulfprdy = '1') then state := s1903;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1902; end if;
when s1903 => state := s1904; 	--12
	mulfpsclr <= '0';
when s1904 => state := s1905; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1905 => 			--14
	if (addfprdy = '1') then state := s1906;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1905; end if;
when s1906 => state := s1907; 	--15
	addfpsclr <= '0';
when s1907 => state := s1908; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1908 => 			--17
	if (addfprdy = '1') then state := s1909;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1908; end if;
when s1909 => state := s1910; 	--18
	addfpsclr <= '0';
when s1910 => state := s1911; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1911 => 			--20
	if (addfprdy = '1') then state := s1912;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1911; end if;
when s1912 => state := s1913; 	--21
	addfpsclr <= '0';
when s1913 => state := s1914; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (142, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1914 => state := s1915; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (222, 12)); -- offset LSB 174
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s1915 => state := s1916;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (223, 12)); -- offset MSB 175
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1916 => state := s1917; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1917 => 			--4
	if (fixed2floatrdy = '1') then state := s1918;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1917; end if;
when s1918 => state := s1919; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1919 => 			--6
	if (mulfprdy = '1') then state := s1920;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1919; end if;
when s1920 => state := s1921; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1921 => 			--8
	if (mulfprdy = '1') then state := s1922;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1921; end if;
when s1922 => state := s1923; 	--9
	mulfpsclr <= '0';
when s1923 => state := s1924; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1924 => 			--11
	if (mulfprdy = '1') then state := s1925;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1924; end if;
when s1925 => state := s1926; 	--12
	mulfpsclr <= '0';
when s1926 => state := s1927; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1927 => 			--14
	if (addfprdy = '1') then state := s1928;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1927; end if;
when s1928 => state := s1929; 	--15
	addfpsclr <= '0';
when s1929 => state := s1930; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1930 => 			--17
	if (addfprdy = '1') then state := s1931;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1930; end if;
when s1931 => state := s1932; 	--18
	addfpsclr <= '0';
when s1932 => state := s1933; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1933 => 			--20
	if (addfprdy = '1') then state := s1934;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1933; end if;
when s1934 => state := s1935; 	--21
	addfpsclr <= '0';
when s1935 => state := s1936; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (143, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1936 => state := s1937; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (224, 12)); -- offset LSB 176
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s1937 => state := s1938;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (225, 12)); -- offset MSB 177
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1938 => state := s1939; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1939 => 			--4
	if (fixed2floatrdy = '1') then state := s1940;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1939; end if;
when s1940 => state := s1941; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1941 => 			--6
	if (mulfprdy = '1') then state := s1942;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1941; end if;
when s1942 => state := s1943; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1943 => 			--8
	if (mulfprdy = '1') then state := s1944;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1943; end if;
when s1944 => state := s1945; 	--9
	mulfpsclr <= '0';
when s1945 => state := s1946; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1946 => 			--11
	if (mulfprdy = '1') then state := s1947;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1946; end if;
when s1947 => state := s1948; 	--12
	mulfpsclr <= '0';
when s1948 => state := s1949; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1949 => 			--14
	if (addfprdy = '1') then state := s1950;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1949; end if;
when s1950 => state := s1951; 	--15
	addfpsclr <= '0';
when s1951 => state := s1952; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1952 => 			--17
	if (addfprdy = '1') then state := s1953;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1952; end if;
when s1953 => state := s1954; 	--18
	addfpsclr <= '0';
when s1954 => state := s1955; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1955 => 			--20
	if (addfprdy = '1') then state := s1956;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1955; end if;
when s1956 => state := s1957; 	--21
	addfpsclr <= '0';
when s1957 => state := s1958; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (144, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1958 => state := s1959; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (226, 12)); -- offset LSB 178
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s1959 => state := s1960;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (227, 12)); -- offset MSB 179
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1960 => state := s1961; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1961 => 			--4
	if (fixed2floatrdy = '1') then state := s1962;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1961; end if;
when s1962 => state := s1963; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1963 => 			--6
	if (mulfprdy = '1') then state := s1964;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1963; end if;
when s1964 => state := s1965; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1965 => 			--8
	if (mulfprdy = '1') then state := s1966;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1965; end if;
when s1966 => state := s1967; 	--9
	mulfpsclr <= '0';
when s1967 => state := s1968; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1968 => 			--11
	if (mulfprdy = '1') then state := s1969;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1968; end if;
when s1969 => state := s1970; 	--12
	mulfpsclr <= '0';
when s1970 => state := s1971; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1971 => 			--14
	if (addfprdy = '1') then state := s1972;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1971; end if;
when s1972 => state := s1973; 	--15
	addfpsclr <= '0';
when s1973 => state := s1974; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1974 => 			--17
	if (addfprdy = '1') then state := s1975;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1974; end if;
when s1975 => state := s1976; 	--18
	addfpsclr <= '0';
when s1976 => state := s1977; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1977 => 			--20
	if (addfprdy = '1') then state := s1978;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1977; end if;
when s1978 => state := s1979; 	--21
	addfpsclr <= '0';
when s1979 => state := s1980; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (145, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s1980 => state := s1981; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (228, 12)); -- offset LSB 180
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s1981 => state := s1982;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (229, 12)); -- offset MSB 181
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s1982 => state := s1983; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s1983 => 			--4
	if (fixed2floatrdy = '1') then state := s1984;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s1983; end if;
when s1984 => state := s1985; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s1985 => 			--6
	if (mulfprdy = '1') then state := s1986;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1985; end if;
when s1986 => state := s1987; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s1987 => 			--8
	if (mulfprdy = '1') then state := s1988;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1987; end if;
when s1988 => state := s1989; 	--9
	mulfpsclr <= '0';
when s1989 => state := s1990; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s1990 => 			--11
	if (mulfprdy = '1') then state := s1991;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s1990; end if;
when s1991 => state := s1992; 	--12
	mulfpsclr <= '0';
when s1992 => state := s1993; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s1993 => 			--14
	if (addfprdy = '1') then state := s1994;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1993; end if;
when s1994 => state := s1995; 	--15
	addfpsclr <= '0';
when s1995 => state := s1996; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s1996 => 			--17
	if (addfprdy = '1') then state := s1997;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1996; end if;
when s1997 => state := s1998; 	--18
	addfpsclr <= '0';
when s1998 => state := s1999; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s1999 => 			--20
	if (addfprdy = '1') then state := s2000;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s1999; end if;
when s2000 => state := s2001; 	--21
	addfpsclr <= '0';
when s2001 => state := s2002; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (146, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2002 => state := s2003; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (230, 12)); -- offset LSB 182
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s2003 => state := s2004;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (231, 12)); -- offset MSB 183
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2004 => state := s2005; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2005 => 			--4
	if (fixed2floatrdy = '1') then state := s2006;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2005; end if;
when s2006 => state := s2007; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2007 => 			--6
	if (mulfprdy = '1') then state := s2008;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2007; end if;
when s2008 => state := s2009; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2009 => 			--8
	if (mulfprdy = '1') then state := s2010;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2009; end if;
when s2010 => state := s2011; 	--9
	mulfpsclr <= '0';
when s2011 => state := s2012; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2012 => 			--11
	if (mulfprdy = '1') then state := s2013;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2012; end if;
when s2013 => state := s2014; 	--12
	mulfpsclr <= '0';
when s2014 => state := s2015; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2015 => 			--14
	if (addfprdy = '1') then state := s2016;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2015; end if;
when s2016 => state := s2017; 	--15
	addfpsclr <= '0';
when s2017 => state := s2018; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2018 => 			--17
	if (addfprdy = '1') then state := s2019;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2018; end if;
when s2019 => state := s2020; 	--18
	addfpsclr <= '0';
when s2020 => state := s2021; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2021 => 			--20
	if (addfprdy = '1') then state := s2022;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2021; end if;
when s2022 => state := s2023; 	--21
	addfpsclr <= '0';
when s2023 => state := s2024; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (147, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2024 => state := s2025; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (232, 12)); -- offset LSB 184
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s2025 => state := s2026;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (233, 12)); -- offset MSB 185
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2026 => state := s2027; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2027 => 			--4
	if (fixed2floatrdy = '1') then state := s2028;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2027; end if;
when s2028 => state := s2029; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2029 => 			--6
	if (mulfprdy = '1') then state := s2030;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2029; end if;
when s2030 => state := s2031; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2031 => 			--8
	if (mulfprdy = '1') then state := s2032;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2031; end if;
when s2032 => state := s2033; 	--9
	mulfpsclr <= '0';
when s2033 => state := s2034; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2034 => 			--11
	if (mulfprdy = '1') then state := s2035;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2034; end if;
when s2035 => state := s2036; 	--12
	mulfpsclr <= '0';
when s2036 => state := s2037; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2037 => 			--14
	if (addfprdy = '1') then state := s2038;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2037; end if;
when s2038 => state := s2039; 	--15
	addfpsclr <= '0';
when s2039 => state := s2040; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2040 => 			--17
	if (addfprdy = '1') then state := s2041;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2040; end if;
when s2041 => state := s2042; 	--18
	addfpsclr <= '0';
when s2042 => state := s2043; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2043 => 			--20
	if (addfprdy = '1') then state := s2044;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2043; end if;
when s2044 => state := s2045; 	--21
	addfpsclr <= '0';
when s2045 => state := s2046; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (148, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2046 => state := s2047; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (234, 12)); -- offset LSB 186
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s2047 => state := s2048;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (235, 12)); -- offset MSB 187
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2048 => state := s2049; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2049 => 			--4
	if (fixed2floatrdy = '1') then state := s2050;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2049; end if;
when s2050 => state := s2051; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2051 => 			--6
	if (mulfprdy = '1') then state := s2052;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2051; end if;
when s2052 => state := s2053; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2053 => 			--8
	if (mulfprdy = '1') then state := s2054;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2053; end if;
when s2054 => state := s2055; 	--9
	mulfpsclr <= '0';
when s2055 => state := s2056; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2056 => 			--11
	if (mulfprdy = '1') then state := s2057;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2056; end if;
when s2057 => state := s2058; 	--12
	mulfpsclr <= '0';
when s2058 => state := s2059; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2059 => 			--14
	if (addfprdy = '1') then state := s2060;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2059; end if;
when s2060 => state := s2061; 	--15
	addfpsclr <= '0';
when s2061 => state := s2062; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2062 => 			--17
	if (addfprdy = '1') then state := s2063;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2062; end if;
when s2063 => state := s2064; 	--18
	addfpsclr <= '0';
when s2064 => state := s2065; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2065 => 			--20
	if (addfprdy = '1') then state := s2066;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2065; end if;
when s2066 => state := s2067; 	--21
	addfpsclr <= '0';
when s2067 => state := s2068; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (149, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2068 => state := s2069; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (236, 12)); -- offset LSB 188
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s2069 => state := s2070;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (237, 12)); -- offset MSB 189
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2070 => state := s2071; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2071 => 			--4
	if (fixed2floatrdy = '1') then state := s2072;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2071; end if;
when s2072 => state := s2073; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2073 => 			--6
	if (mulfprdy = '1') then state := s2074;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2073; end if;
when s2074 => state := s2075; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2075 => 			--8
	if (mulfprdy = '1') then state := s2076;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2075; end if;
when s2076 => state := s2077; 	--9
	mulfpsclr <= '0';
when s2077 => state := s2078; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2078 => 			--11
	if (mulfprdy = '1') then state := s2079;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2078; end if;
when s2079 => state := s2080; 	--12
	mulfpsclr <= '0';
when s2080 => state := s2081; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2081 => 			--14
	if (addfprdy = '1') then state := s2082;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2081; end if;
when s2082 => state := s2083; 	--15
	addfpsclr <= '0';
when s2083 => state := s2084; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2084 => 			--17
	if (addfprdy = '1') then state := s2085;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2084; end if;
when s2085 => state := s2086; 	--18
	addfpsclr <= '0';
when s2086 => state := s2087; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2087 => 			--20
	if (addfprdy = '1') then state := s2088;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2087; end if;
when s2088 => state := s2089; 	--21
	addfpsclr <= '0';
when s2089 => state := s2090; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (150, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2090 => state := s2091; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (238, 12)); -- offset LSB 190
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s2091 => state := s2092;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (239, 12)); -- offset MSB 191
	addra <= std_logic_vector (to_unsigned (2, 10)); -- OCCrowI 2
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2092 => state := s2093; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2093 => 			--4
	if (fixed2floatrdy = '1') then state := s2094;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2093; end if;
when s2094 => state := s2095; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2095 => 			--6
	if (mulfprdy = '1') then state := s2096;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2095; end if;
when s2096 => state := s2097; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2097 => 			--8
	if (mulfprdy = '1') then state := s2098;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2097; end if;
when s2098 => state := s2099; 	--9
	mulfpsclr <= '0';
when s2099 => state := s2100; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2100 => 			--11
	if (mulfprdy = '1') then state := s2101;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2100; end if;
when s2101 => state := s2102; 	--12
	mulfpsclr <= '0';
when s2102 => state := s2103; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2103 => 			--14
	if (addfprdy = '1') then state := s2104;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2103; end if;
when s2104 => state := s2105; 	--15
	addfpsclr <= '0';
when s2105 => state := s2106; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2106 => 			--17
	if (addfprdy = '1') then state := s2107;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2106; end if;
when s2107 => state := s2108; 	--18
	addfpsclr <= '0';
when s2108 => state := s2109; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2109 => 			--20
	if (addfprdy = '1') then state := s2110;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2109; end if;
when s2110 => state := s2111; 	--21
	addfpsclr <= '0';
when s2111 => state := s2112; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (151, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2112 => state := s2113; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (240, 12)); -- offset LSB 192
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s2113 => state := s2114;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (241, 12)); -- offset MSB 193
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2114 => state := s2115; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2115 => 			--4
	if (fixed2floatrdy = '1') then state := s2116;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2115; end if;
when s2116 => state := s2117; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2117 => 			--6
	if (mulfprdy = '1') then state := s2118;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2117; end if;
when s2118 => state := s2119; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2119 => 			--8
	if (mulfprdy = '1') then state := s2120;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2119; end if;
when s2120 => state := s2121; 	--9
	mulfpsclr <= '0';
when s2121 => state := s2122; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2122 => 			--11
	if (mulfprdy = '1') then state := s2123;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2122; end if;
when s2123 => state := s2124; 	--12
	mulfpsclr <= '0';
when s2124 => state := s2125; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2125 => 			--14
	if (addfprdy = '1') then state := s2126;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2125; end if;
when s2126 => state := s2127; 	--15
	addfpsclr <= '0';
when s2127 => state := s2128; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2128 => 			--17
	if (addfprdy = '1') then state := s2129;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2128; end if;
when s2129 => state := s2130; 	--18
	addfpsclr <= '0';
when s2130 => state := s2131; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2131 => 			--20
	if (addfprdy = '1') then state := s2132;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2131; end if;
when s2132 => state := s2133; 	--21
	addfpsclr <= '0';
when s2133 => state := s2134; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (152, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2134 => state := s2135; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (242, 12)); -- offset LSB 194
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s2135 => state := s2136;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (243, 12)); -- offset MSB 195
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2136 => state := s2137; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2137 => 			--4
	if (fixed2floatrdy = '1') then state := s2138;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2137; end if;
when s2138 => state := s2139; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2139 => 			--6
	if (mulfprdy = '1') then state := s2140;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2139; end if;
when s2140 => state := s2141; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2141 => 			--8
	if (mulfprdy = '1') then state := s2142;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2141; end if;
when s2142 => state := s2143; 	--9
	mulfpsclr <= '0';
when s2143 => state := s2144; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2144 => 			--11
	if (mulfprdy = '1') then state := s2145;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2144; end if;
when s2145 => state := s2146; 	--12
	mulfpsclr <= '0';
when s2146 => state := s2147; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2147 => 			--14
	if (addfprdy = '1') then state := s2148;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2147; end if;
when s2148 => state := s2149; 	--15
	addfpsclr <= '0';
when s2149 => state := s2150; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2150 => 			--17
	if (addfprdy = '1') then state := s2151;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2150; end if;
when s2151 => state := s2152; 	--18
	addfpsclr <= '0';
when s2152 => state := s2153; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2153 => 			--20
	if (addfprdy = '1') then state := s2154;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2153; end if;
when s2154 => state := s2155; 	--21
	addfpsclr <= '0';
when s2155 => state := s2156; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (153, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2156 => state := s2157; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (244, 12)); -- offset LSB 196
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s2157 => state := s2158;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (245, 12)); -- offset MSB 197
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2158 => state := s2159; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2159 => 			--4
	if (fixed2floatrdy = '1') then state := s2160;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2159; end if;
when s2160 => state := s2161; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2161 => 			--6
	if (mulfprdy = '1') then state := s2162;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2161; end if;
when s2162 => state := s2163; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2163 => 			--8
	if (mulfprdy = '1') then state := s2164;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2163; end if;
when s2164 => state := s2165; 	--9
	mulfpsclr <= '0';
when s2165 => state := s2166; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2166 => 			--11
	if (mulfprdy = '1') then state := s2167;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2166; end if;
when s2167 => state := s2168; 	--12
	mulfpsclr <= '0';
when s2168 => state := s2169; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2169 => 			--14
	if (addfprdy = '1') then state := s2170;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2169; end if;
when s2170 => state := s2171; 	--15
	addfpsclr <= '0';
when s2171 => state := s2172; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2172 => 			--17
	if (addfprdy = '1') then state := s2173;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2172; end if;
when s2173 => state := s2174; 	--18
	addfpsclr <= '0';
when s2174 => state := s2175; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2175 => 			--20
	if (addfprdy = '1') then state := s2176;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2175; end if;
when s2176 => state := s2177; 	--21
	addfpsclr <= '0';
when s2177 => state := s2178; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (154, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2178 => state := s2179; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (246, 12)); -- offset LSB 198
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s2179 => state := s2180;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (247, 12)); -- offset MSB 199
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2180 => state := s2181; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2181 => 			--4
	if (fixed2floatrdy = '1') then state := s2182;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2181; end if;
when s2182 => state := s2183; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2183 => 			--6
	if (mulfprdy = '1') then state := s2184;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2183; end if;
when s2184 => state := s2185; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2185 => 			--8
	if (mulfprdy = '1') then state := s2186;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2185; end if;
when s2186 => state := s2187; 	--9
	mulfpsclr <= '0';
when s2187 => state := s2188; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2188 => 			--11
	if (mulfprdy = '1') then state := s2189;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2188; end if;
when s2189 => state := s2190; 	--12
	mulfpsclr <= '0';
when s2190 => state := s2191; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2191 => 			--14
	if (addfprdy = '1') then state := s2192;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2191; end if;
when s2192 => state := s2193; 	--15
	addfpsclr <= '0';
when s2193 => state := s2194; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2194 => 			--17
	if (addfprdy = '1') then state := s2195;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2194; end if;
when s2195 => state := s2196; 	--18
	addfpsclr <= '0';
when s2196 => state := s2197; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2197 => 			--20
	if (addfprdy = '1') then state := s2198;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2197; end if;
when s2198 => state := s2199; 	--21
	addfpsclr <= '0';
when s2199 => state := s2200; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (155, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2200 => state := s2201; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (248, 12)); -- offset LSB 200
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s2201 => state := s2202;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (249, 12)); -- offset MSB 201
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2202 => state := s2203; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2203 => 			--4
	if (fixed2floatrdy = '1') then state := s2204;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2203; end if;
when s2204 => state := s2205; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2205 => 			--6
	if (mulfprdy = '1') then state := s2206;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2205; end if;
when s2206 => state := s2207; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2207 => 			--8
	if (mulfprdy = '1') then state := s2208;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2207; end if;
when s2208 => state := s2209; 	--9
	mulfpsclr <= '0';
when s2209 => state := s2210; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2210 => 			--11
	if (mulfprdy = '1') then state := s2211;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2210; end if;
when s2211 => state := s2212; 	--12
	mulfpsclr <= '0';
when s2212 => state := s2213; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2213 => 			--14
	if (addfprdy = '1') then state := s2214;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2213; end if;
when s2214 => state := s2215; 	--15
	addfpsclr <= '0';
when s2215 => state := s2216; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2216 => 			--17
	if (addfprdy = '1') then state := s2217;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2216; end if;
when s2217 => state := s2218; 	--18
	addfpsclr <= '0';
when s2218 => state := s2219; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2219 => 			--20
	if (addfprdy = '1') then state := s2220;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2219; end if;
when s2220 => state := s2221; 	--21
	addfpsclr <= '0';
when s2221 => state := s2222; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (156, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2222 => state := s2223; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (250, 12)); -- offset LSB 202
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s2223 => state := s2224;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (251, 12)); -- offset MSB 203
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2224 => state := s2225; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2225 => 			--4
	if (fixed2floatrdy = '1') then state := s2226;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2225; end if;
when s2226 => state := s2227; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2227 => 			--6
	if (mulfprdy = '1') then state := s2228;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2227; end if;
when s2228 => state := s2229; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2229 => 			--8
	if (mulfprdy = '1') then state := s2230;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2229; end if;
when s2230 => state := s2231; 	--9
	mulfpsclr <= '0';
when s2231 => state := s2232; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2232 => 			--11
	if (mulfprdy = '1') then state := s2233;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2232; end if;
when s2233 => state := s2234; 	--12
	mulfpsclr <= '0';
when s2234 => state := s2235; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2235 => 			--14
	if (addfprdy = '1') then state := s2236;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2235; end if;
when s2236 => state := s2237; 	--15
	addfpsclr <= '0';
when s2237 => state := s2238; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2238 => 			--17
	if (addfprdy = '1') then state := s2239;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2238; end if;
when s2239 => state := s2240; 	--18
	addfpsclr <= '0';
when s2240 => state := s2241; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2241 => 			--20
	if (addfprdy = '1') then state := s2242;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2241; end if;
when s2242 => state := s2243; 	--21
	addfpsclr <= '0';
when s2243 => state := s2244; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (157, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2244 => state := s2245; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (252, 12)); -- offset LSB 204
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s2245 => state := s2246;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (253, 12)); -- offset MSB 205
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2246 => state := s2247; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2247 => 			--4
	if (fixed2floatrdy = '1') then state := s2248;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2247; end if;
when s2248 => state := s2249; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2249 => 			--6
	if (mulfprdy = '1') then state := s2250;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2249; end if;
when s2250 => state := s2251; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2251 => 			--8
	if (mulfprdy = '1') then state := s2252;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2251; end if;
when s2252 => state := s2253; 	--9
	mulfpsclr <= '0';
when s2253 => state := s2254; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2254 => 			--11
	if (mulfprdy = '1') then state := s2255;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2254; end if;
when s2255 => state := s2256; 	--12
	mulfpsclr <= '0';
when s2256 => state := s2257; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2257 => 			--14
	if (addfprdy = '1') then state := s2258;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2257; end if;
when s2258 => state := s2259; 	--15
	addfpsclr <= '0';
when s2259 => state := s2260; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2260 => 			--17
	if (addfprdy = '1') then state := s2261;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2260; end if;
when s2261 => state := s2262; 	--18
	addfpsclr <= '0';
when s2262 => state := s2263; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2263 => 			--20
	if (addfprdy = '1') then state := s2264;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2263; end if;
when s2264 => state := s2265; 	--21
	addfpsclr <= '0';
when s2265 => state := s2266; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (158, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2266 => state := s2267; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (254, 12)); -- offset LSB 206
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s2267 => state := s2268;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (255, 12)); -- offset MSB 207
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2268 => state := s2269; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2269 => 			--4
	if (fixed2floatrdy = '1') then state := s2270;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2269; end if;
when s2270 => state := s2271; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2271 => 			--6
	if (mulfprdy = '1') then state := s2272;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2271; end if;
when s2272 => state := s2273; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2273 => 			--8
	if (mulfprdy = '1') then state := s2274;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2273; end if;
when s2274 => state := s2275; 	--9
	mulfpsclr <= '0';
when s2275 => state := s2276; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2276 => 			--11
	if (mulfprdy = '1') then state := s2277;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2276; end if;
when s2277 => state := s2278; 	--12
	mulfpsclr <= '0';
when s2278 => state := s2279; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2279 => 			--14
	if (addfprdy = '1') then state := s2280;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2279; end if;
when s2280 => state := s2281; 	--15
	addfpsclr <= '0';
when s2281 => state := s2282; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2282 => 			--17
	if (addfprdy = '1') then state := s2283;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2282; end if;
when s2283 => state := s2284; 	--18
	addfpsclr <= '0';
when s2284 => state := s2285; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2285 => 			--20
	if (addfprdy = '1') then state := s2286;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2285; end if;
when s2286 => state := s2287; 	--21
	addfpsclr <= '0';
when s2287 => state := s2288; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (159, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2288 => state := s2289; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (256, 12)); -- offset LSB 208
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s2289 => state := s2290;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (257, 12)); -- offset MSB 209
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2290 => state := s2291; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2291 => 			--4
	if (fixed2floatrdy = '1') then state := s2292;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2291; end if;
when s2292 => state := s2293; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2293 => 			--6
	if (mulfprdy = '1') then state := s2294;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2293; end if;
when s2294 => state := s2295; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2295 => 			--8
	if (mulfprdy = '1') then state := s2296;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2295; end if;
when s2296 => state := s2297; 	--9
	mulfpsclr <= '0';
when s2297 => state := s2298; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2298 => 			--11
	if (mulfprdy = '1') then state := s2299;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2298; end if;
when s2299 => state := s2300; 	--12
	mulfpsclr <= '0';
when s2300 => state := s2301; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2301 => 			--14
	if (addfprdy = '1') then state := s2302;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2301; end if;
when s2302 => state := s2303; 	--15
	addfpsclr <= '0';
when s2303 => state := s2304; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2304 => 			--17
	if (addfprdy = '1') then state := s2305;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2304; end if;
when s2305 => state := s2306; 	--18
	addfpsclr <= '0';
when s2306 => state := s2307; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2307 => 			--20
	if (addfprdy = '1') then state := s2308;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2307; end if;
when s2308 => state := s2309; 	--21
	addfpsclr <= '0';
when s2309 => state := s2310; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (160, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2310 => state := s2311; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (258, 12)); -- offset LSB 210
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s2311 => state := s2312;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (259, 12)); -- offset MSB 211
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2312 => state := s2313; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2313 => 			--4
	if (fixed2floatrdy = '1') then state := s2314;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2313; end if;
when s2314 => state := s2315; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2315 => 			--6
	if (mulfprdy = '1') then state := s2316;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2315; end if;
when s2316 => state := s2317; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2317 => 			--8
	if (mulfprdy = '1') then state := s2318;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2317; end if;
when s2318 => state := s2319; 	--9
	mulfpsclr <= '0';
when s2319 => state := s2320; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2320 => 			--11
	if (mulfprdy = '1') then state := s2321;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2320; end if;
when s2321 => state := s2322; 	--12
	mulfpsclr <= '0';
when s2322 => state := s2323; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2323 => 			--14
	if (addfprdy = '1') then state := s2324;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2323; end if;
when s2324 => state := s2325; 	--15
	addfpsclr <= '0';
when s2325 => state := s2326; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2326 => 			--17
	if (addfprdy = '1') then state := s2327;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2326; end if;
when s2327 => state := s2328; 	--18
	addfpsclr <= '0';
when s2328 => state := s2329; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2329 => 			--20
	if (addfprdy = '1') then state := s2330;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2329; end if;
when s2330 => state := s2331; 	--21
	addfpsclr <= '0';
when s2331 => state := s2332; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (161, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2332 => state := s2333; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (260, 12)); -- offset LSB 212
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s2333 => state := s2334;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (261, 12)); -- offset MSB 213
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2334 => state := s2335; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2335 => 			--4
	if (fixed2floatrdy = '1') then state := s2336;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2335; end if;
when s2336 => state := s2337; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2337 => 			--6
	if (mulfprdy = '1') then state := s2338;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2337; end if;
when s2338 => state := s2339; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2339 => 			--8
	if (mulfprdy = '1') then state := s2340;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2339; end if;
when s2340 => state := s2341; 	--9
	mulfpsclr <= '0';
when s2341 => state := s2342; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2342 => 			--11
	if (mulfprdy = '1') then state := s2343;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2342; end if;
when s2343 => state := s2344; 	--12
	mulfpsclr <= '0';
when s2344 => state := s2345; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2345 => 			--14
	if (addfprdy = '1') then state := s2346;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2345; end if;
when s2346 => state := s2347; 	--15
	addfpsclr <= '0';
when s2347 => state := s2348; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2348 => 			--17
	if (addfprdy = '1') then state := s2349;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2348; end if;
when s2349 => state := s2350; 	--18
	addfpsclr <= '0';
when s2350 => state := s2351; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2351 => 			--20
	if (addfprdy = '1') then state := s2352;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2351; end if;
when s2352 => state := s2353; 	--21
	addfpsclr <= '0';
when s2353 => state := s2354; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (162, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2354 => state := s2355; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (262, 12)); -- offset LSB 214
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s2355 => state := s2356;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (263, 12)); -- offset MSB 215
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2356 => state := s2357; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2357 => 			--4
	if (fixed2floatrdy = '1') then state := s2358;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2357; end if;
when s2358 => state := s2359; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2359 => 			--6
	if (mulfprdy = '1') then state := s2360;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2359; end if;
when s2360 => state := s2361; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2361 => 			--8
	if (mulfprdy = '1') then state := s2362;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2361; end if;
when s2362 => state := s2363; 	--9
	mulfpsclr <= '0';
when s2363 => state := s2364; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2364 => 			--11
	if (mulfprdy = '1') then state := s2365;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2364; end if;
when s2365 => state := s2366; 	--12
	mulfpsclr <= '0';
when s2366 => state := s2367; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2367 => 			--14
	if (addfprdy = '1') then state := s2368;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2367; end if;
when s2368 => state := s2369; 	--15
	addfpsclr <= '0';
when s2369 => state := s2370; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2370 => 			--17
	if (addfprdy = '1') then state := s2371;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2370; end if;
when s2371 => state := s2372; 	--18
	addfpsclr <= '0';
when s2372 => state := s2373; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2373 => 			--20
	if (addfprdy = '1') then state := s2374;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2373; end if;
when s2374 => state := s2375; 	--21
	addfpsclr <= '0';
when s2375 => state := s2376; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (163, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2376 => state := s2377; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (264, 12)); -- offset LSB 216
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s2377 => state := s2378;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (265, 12)); -- offset MSB 217
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2378 => state := s2379; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2379 => 			--4
	if (fixed2floatrdy = '1') then state := s2380;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2379; end if;
when s2380 => state := s2381; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2381 => 			--6
	if (mulfprdy = '1') then state := s2382;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2381; end if;
when s2382 => state := s2383; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2383 => 			--8
	if (mulfprdy = '1') then state := s2384;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2383; end if;
when s2384 => state := s2385; 	--9
	mulfpsclr <= '0';
when s2385 => state := s2386; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2386 => 			--11
	if (mulfprdy = '1') then state := s2387;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2386; end if;
when s2387 => state := s2388; 	--12
	mulfpsclr <= '0';
when s2388 => state := s2389; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2389 => 			--14
	if (addfprdy = '1') then state := s2390;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2389; end if;
when s2390 => state := s2391; 	--15
	addfpsclr <= '0';
when s2391 => state := s2392; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2392 => 			--17
	if (addfprdy = '1') then state := s2393;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2392; end if;
when s2393 => state := s2394; 	--18
	addfpsclr <= '0';
when s2394 => state := s2395; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2395 => 			--20
	if (addfprdy = '1') then state := s2396;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2395; end if;
when s2396 => state := s2397; 	--21
	addfpsclr <= '0';
when s2397 => state := s2398; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (164, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2398 => state := s2399; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (266, 12)); -- offset LSB 218
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s2399 => state := s2400;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (267, 12)); -- offset MSB 219
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2400 => state := s2401; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2401 => 			--4
	if (fixed2floatrdy = '1') then state := s2402;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2401; end if;
when s2402 => state := s2403; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2403 => 			--6
	if (mulfprdy = '1') then state := s2404;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2403; end if;
when s2404 => state := s2405; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2405 => 			--8
	if (mulfprdy = '1') then state := s2406;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2405; end if;
when s2406 => state := s2407; 	--9
	mulfpsclr <= '0';
when s2407 => state := s2408; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2408 => 			--11
	if (mulfprdy = '1') then state := s2409;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2408; end if;
when s2409 => state := s2410; 	--12
	mulfpsclr <= '0';
when s2410 => state := s2411; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2411 => 			--14
	if (addfprdy = '1') then state := s2412;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2411; end if;
when s2412 => state := s2413; 	--15
	addfpsclr <= '0';
when s2413 => state := s2414; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2414 => 			--17
	if (addfprdy = '1') then state := s2415;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2414; end if;
when s2415 => state := s2416; 	--18
	addfpsclr <= '0';
when s2416 => state := s2417; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2417 => 			--20
	if (addfprdy = '1') then state := s2418;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2417; end if;
when s2418 => state := s2419; 	--21
	addfpsclr <= '0';
when s2419 => state := s2420; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (165, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2420 => state := s2421; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (268, 12)); -- offset LSB 220
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s2421 => state := s2422;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (269, 12)); -- offset MSB 221
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2422 => state := s2423; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2423 => 			--4
	if (fixed2floatrdy = '1') then state := s2424;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2423; end if;
when s2424 => state := s2425; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2425 => 			--6
	if (mulfprdy = '1') then state := s2426;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2425; end if;
when s2426 => state := s2427; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2427 => 			--8
	if (mulfprdy = '1') then state := s2428;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2427; end if;
when s2428 => state := s2429; 	--9
	mulfpsclr <= '0';
when s2429 => state := s2430; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2430 => 			--11
	if (mulfprdy = '1') then state := s2431;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2430; end if;
when s2431 => state := s2432; 	--12
	mulfpsclr <= '0';
when s2432 => state := s2433; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2433 => 			--14
	if (addfprdy = '1') then state := s2434;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2433; end if;
when s2434 => state := s2435; 	--15
	addfpsclr <= '0';
when s2435 => state := s2436; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2436 => 			--17
	if (addfprdy = '1') then state := s2437;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2436; end if;
when s2437 => state := s2438; 	--18
	addfpsclr <= '0';
when s2438 => state := s2439; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2439 => 			--20
	if (addfprdy = '1') then state := s2440;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2439; end if;
when s2440 => state := s2441; 	--21
	addfpsclr <= '0';
when s2441 => state := s2442; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (166, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2442 => state := s2443; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (270, 12)); -- offset LSB 222
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s2443 => state := s2444;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (271, 12)); -- offset MSB 223
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2444 => state := s2445; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2445 => 			--4
	if (fixed2floatrdy = '1') then state := s2446;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2445; end if;
when s2446 => state := s2447; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2447 => 			--6
	if (mulfprdy = '1') then state := s2448;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2447; end if;
when s2448 => state := s2449; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2449 => 			--8
	if (mulfprdy = '1') then state := s2450;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2449; end if;
when s2450 => state := s2451; 	--9
	mulfpsclr <= '0';
when s2451 => state := s2452; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2452 => 			--11
	if (mulfprdy = '1') then state := s2453;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2452; end if;
when s2453 => state := s2454; 	--12
	mulfpsclr <= '0';
when s2454 => state := s2455; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2455 => 			--14
	if (addfprdy = '1') then state := s2456;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2455; end if;
when s2456 => state := s2457; 	--15
	addfpsclr <= '0';
when s2457 => state := s2458; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2458 => 			--17
	if (addfprdy = '1') then state := s2459;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2458; end if;
when s2459 => state := s2460; 	--18
	addfpsclr <= '0';
when s2460 => state := s2461; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2461 => 			--20
	if (addfprdy = '1') then state := s2462;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2461; end if;
when s2462 => state := s2463; 	--21
	addfpsclr <= '0';
when s2463 => state := s2464; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (167, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2464 => state := s2465; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (272, 12)); -- offset LSB 224
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s2465 => state := s2466;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (273, 12)); -- offset MSB 225
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2466 => state := s2467; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2467 => 			--4
	if (fixed2floatrdy = '1') then state := s2468;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2467; end if;
when s2468 => state := s2469; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2469 => 			--6
	if (mulfprdy = '1') then state := s2470;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2469; end if;
when s2470 => state := s2471; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2471 => 			--8
	if (mulfprdy = '1') then state := s2472;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2471; end if;
when s2472 => state := s2473; 	--9
	mulfpsclr <= '0';
when s2473 => state := s2474; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2474 => 			--11
	if (mulfprdy = '1') then state := s2475;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2474; end if;
when s2475 => state := s2476; 	--12
	mulfpsclr <= '0';
when s2476 => state := s2477; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2477 => 			--14
	if (addfprdy = '1') then state := s2478;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2477; end if;
when s2478 => state := s2479; 	--15
	addfpsclr <= '0';
when s2479 => state := s2480; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2480 => 			--17
	if (addfprdy = '1') then state := s2481;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2480; end if;
when s2481 => state := s2482; 	--18
	addfpsclr <= '0';
when s2482 => state := s2483; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2483 => 			--20
	if (addfprdy = '1') then state := s2484;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2483; end if;
when s2484 => state := s2485; 	--21
	addfpsclr <= '0';
when s2485 => state := s2486; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (168, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2486 => state := s2487; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (274, 12)); -- offset LSB 226
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s2487 => state := s2488;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (275, 12)); -- offset MSB 227
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2488 => state := s2489; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2489 => 			--4
	if (fixed2floatrdy = '1') then state := s2490;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2489; end if;
when s2490 => state := s2491; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2491 => 			--6
	if (mulfprdy = '1') then state := s2492;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2491; end if;
when s2492 => state := s2493; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2493 => 			--8
	if (mulfprdy = '1') then state := s2494;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2493; end if;
when s2494 => state := s2495; 	--9
	mulfpsclr <= '0';
when s2495 => state := s2496; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2496 => 			--11
	if (mulfprdy = '1') then state := s2497;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2496; end if;
when s2497 => state := s2498; 	--12
	mulfpsclr <= '0';
when s2498 => state := s2499; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2499 => 			--14
	if (addfprdy = '1') then state := s2500;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2499; end if;
when s2500 => state := s2501; 	--15
	addfpsclr <= '0';
when s2501 => state := s2502; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2502 => 			--17
	if (addfprdy = '1') then state := s2503;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2502; end if;
when s2503 => state := s2504; 	--18
	addfpsclr <= '0';
when s2504 => state := s2505; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2505 => 			--20
	if (addfprdy = '1') then state := s2506;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2505; end if;
when s2506 => state := s2507; 	--21
	addfpsclr <= '0';
when s2507 => state := s2508; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (169, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2508 => state := s2509; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (276, 12)); -- offset LSB 228
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s2509 => state := s2510;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (277, 12)); -- offset MSB 229
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2510 => state := s2511; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2511 => 			--4
	if (fixed2floatrdy = '1') then state := s2512;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2511; end if;
when s2512 => state := s2513; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2513 => 			--6
	if (mulfprdy = '1') then state := s2514;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2513; end if;
when s2514 => state := s2515; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2515 => 			--8
	if (mulfprdy = '1') then state := s2516;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2515; end if;
when s2516 => state := s2517; 	--9
	mulfpsclr <= '0';
when s2517 => state := s2518; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2518 => 			--11
	if (mulfprdy = '1') then state := s2519;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2518; end if;
when s2519 => state := s2520; 	--12
	mulfpsclr <= '0';
when s2520 => state := s2521; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2521 => 			--14
	if (addfprdy = '1') then state := s2522;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2521; end if;
when s2522 => state := s2523; 	--15
	addfpsclr <= '0';
when s2523 => state := s2524; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2524 => 			--17
	if (addfprdy = '1') then state := s2525;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2524; end if;
when s2525 => state := s2526; 	--18
	addfpsclr <= '0';
when s2526 => state := s2527; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2527 => 			--20
	if (addfprdy = '1') then state := s2528;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2527; end if;
when s2528 => state := s2529; 	--21
	addfpsclr <= '0';
when s2529 => state := s2530; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (170, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2530 => state := s2531; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (278, 12)); -- offset LSB 230
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s2531 => state := s2532;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (279, 12)); -- offset MSB 231
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2532 => state := s2533; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2533 => 			--4
	if (fixed2floatrdy = '1') then state := s2534;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2533; end if;
when s2534 => state := s2535; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2535 => 			--6
	if (mulfprdy = '1') then state := s2536;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2535; end if;
when s2536 => state := s2537; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2537 => 			--8
	if (mulfprdy = '1') then state := s2538;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2537; end if;
when s2538 => state := s2539; 	--9
	mulfpsclr <= '0';
when s2539 => state := s2540; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2540 => 			--11
	if (mulfprdy = '1') then state := s2541;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2540; end if;
when s2541 => state := s2542; 	--12
	mulfpsclr <= '0';
when s2542 => state := s2543; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2543 => 			--14
	if (addfprdy = '1') then state := s2544;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2543; end if;
when s2544 => state := s2545; 	--15
	addfpsclr <= '0';
when s2545 => state := s2546; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2546 => 			--17
	if (addfprdy = '1') then state := s2547;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2546; end if;
when s2547 => state := s2548; 	--18
	addfpsclr <= '0';
when s2548 => state := s2549; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2549 => 			--20
	if (addfprdy = '1') then state := s2550;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2549; end if;
when s2550 => state := s2551; 	--21
	addfpsclr <= '0';
when s2551 => state := s2552; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (171, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2552 => state := s2553; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (280, 12)); -- offset LSB 232
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s2553 => state := s2554;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (281, 12)); -- offset MSB 233
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2554 => state := s2555; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2555 => 			--4
	if (fixed2floatrdy = '1') then state := s2556;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2555; end if;
when s2556 => state := s2557; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2557 => 			--6
	if (mulfprdy = '1') then state := s2558;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2557; end if;
when s2558 => state := s2559; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2559 => 			--8
	if (mulfprdy = '1') then state := s2560;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2559; end if;
when s2560 => state := s2561; 	--9
	mulfpsclr <= '0';
when s2561 => state := s2562; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2562 => 			--11
	if (mulfprdy = '1') then state := s2563;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2562; end if;
when s2563 => state := s2564; 	--12
	mulfpsclr <= '0';
when s2564 => state := s2565; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2565 => 			--14
	if (addfprdy = '1') then state := s2566;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2565; end if;
when s2566 => state := s2567; 	--15
	addfpsclr <= '0';
when s2567 => state := s2568; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2568 => 			--17
	if (addfprdy = '1') then state := s2569;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2568; end if;
when s2569 => state := s2570; 	--18
	addfpsclr <= '0';
when s2570 => state := s2571; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2571 => 			--20
	if (addfprdy = '1') then state := s2572;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2571; end if;
when s2572 => state := s2573; 	--21
	addfpsclr <= '0';
when s2573 => state := s2574; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (172, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2574 => state := s2575; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (282, 12)); -- offset LSB 234
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s2575 => state := s2576;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (283, 12)); -- offset MSB 235
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2576 => state := s2577; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2577 => 			--4
	if (fixed2floatrdy = '1') then state := s2578;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2577; end if;
when s2578 => state := s2579; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2579 => 			--6
	if (mulfprdy = '1') then state := s2580;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2579; end if;
when s2580 => state := s2581; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2581 => 			--8
	if (mulfprdy = '1') then state := s2582;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2581; end if;
when s2582 => state := s2583; 	--9
	mulfpsclr <= '0';
when s2583 => state := s2584; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2584 => 			--11
	if (mulfprdy = '1') then state := s2585;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2584; end if;
when s2585 => state := s2586; 	--12
	mulfpsclr <= '0';
when s2586 => state := s2587; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2587 => 			--14
	if (addfprdy = '1') then state := s2588;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2587; end if;
when s2588 => state := s2589; 	--15
	addfpsclr <= '0';
when s2589 => state := s2590; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2590 => 			--17
	if (addfprdy = '1') then state := s2591;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2590; end if;
when s2591 => state := s2592; 	--18
	addfpsclr <= '0';
when s2592 => state := s2593; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2593 => 			--20
	if (addfprdy = '1') then state := s2594;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2593; end if;
when s2594 => state := s2595; 	--21
	addfpsclr <= '0';
when s2595 => state := s2596; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (173, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2596 => state := s2597; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (284, 12)); -- offset LSB 236
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s2597 => state := s2598;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (285, 12)); -- offset MSB 237
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2598 => state := s2599; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2599 => 			--4
	if (fixed2floatrdy = '1') then state := s2600;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2599; end if;
when s2600 => state := s2601; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2601 => 			--6
	if (mulfprdy = '1') then state := s2602;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2601; end if;
when s2602 => state := s2603; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2603 => 			--8
	if (mulfprdy = '1') then state := s2604;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2603; end if;
when s2604 => state := s2605; 	--9
	mulfpsclr <= '0';
when s2605 => state := s2606; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2606 => 			--11
	if (mulfprdy = '1') then state := s2607;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2606; end if;
when s2607 => state := s2608; 	--12
	mulfpsclr <= '0';
when s2608 => state := s2609; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2609 => 			--14
	if (addfprdy = '1') then state := s2610;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2609; end if;
when s2610 => state := s2611; 	--15
	addfpsclr <= '0';
when s2611 => state := s2612; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2612 => 			--17
	if (addfprdy = '1') then state := s2613;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2612; end if;
when s2613 => state := s2614; 	--18
	addfpsclr <= '0';
when s2614 => state := s2615; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2615 => 			--20
	if (addfprdy = '1') then state := s2616;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2615; end if;
when s2616 => state := s2617; 	--21
	addfpsclr <= '0';
when s2617 => state := s2618; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (174, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2618 => state := s2619; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (286, 12)); -- offset LSB 238
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s2619 => state := s2620;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (287, 12)); -- offset MSB 239
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2620 => state := s2621; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2621 => 			--4
	if (fixed2floatrdy = '1') then state := s2622;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2621; end if;
when s2622 => state := s2623; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2623 => 			--6
	if (mulfprdy = '1') then state := s2624;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2623; end if;
when s2624 => state := s2625; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2625 => 			--8
	if (mulfprdy = '1') then state := s2626;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2625; end if;
when s2626 => state := s2627; 	--9
	mulfpsclr <= '0';
when s2627 => state := s2628; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2628 => 			--11
	if (mulfprdy = '1') then state := s2629;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2628; end if;
when s2629 => state := s2630; 	--12
	mulfpsclr <= '0';
when s2630 => state := s2631; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2631 => 			--14
	if (addfprdy = '1') then state := s2632;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2631; end if;
when s2632 => state := s2633; 	--15
	addfpsclr <= '0';
when s2633 => state := s2634; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2634 => 			--17
	if (addfprdy = '1') then state := s2635;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2634; end if;
when s2635 => state := s2636; 	--18
	addfpsclr <= '0';
when s2636 => state := s2637; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2637 => 			--20
	if (addfprdy = '1') then state := s2638;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2637; end if;
when s2638 => state := s2639; 	--21
	addfpsclr <= '0';
when s2639 => state := s2640; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (175, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2640 => state := s2641; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (288, 12)); -- offset LSB 240
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s2641 => state := s2642;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (289, 12)); -- offset MSB 241
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2642 => state := s2643; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2643 => 			--4
	if (fixed2floatrdy = '1') then state := s2644;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2643; end if;
when s2644 => state := s2645; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2645 => 			--6
	if (mulfprdy = '1') then state := s2646;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2645; end if;
when s2646 => state := s2647; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2647 => 			--8
	if (mulfprdy = '1') then state := s2648;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2647; end if;
when s2648 => state := s2649; 	--9
	mulfpsclr <= '0';
when s2649 => state := s2650; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2650 => 			--11
	if (mulfprdy = '1') then state := s2651;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2650; end if;
when s2651 => state := s2652; 	--12
	mulfpsclr <= '0';
when s2652 => state := s2653; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2653 => 			--14
	if (addfprdy = '1') then state := s2654;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2653; end if;
when s2654 => state := s2655; 	--15
	addfpsclr <= '0';
when s2655 => state := s2656; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2656 => 			--17
	if (addfprdy = '1') then state := s2657;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2656; end if;
when s2657 => state := s2658; 	--18
	addfpsclr <= '0';
when s2658 => state := s2659; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2659 => 			--20
	if (addfprdy = '1') then state := s2660;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2659; end if;
when s2660 => state := s2661; 	--21
	addfpsclr <= '0';
when s2661 => state := s2662; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (176, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2662 => state := s2663; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (290, 12)); -- offset LSB 242
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s2663 => state := s2664;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (291, 12)); -- offset MSB 243
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2664 => state := s2665; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2665 => 			--4
	if (fixed2floatrdy = '1') then state := s2666;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2665; end if;
when s2666 => state := s2667; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2667 => 			--6
	if (mulfprdy = '1') then state := s2668;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2667; end if;
when s2668 => state := s2669; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2669 => 			--8
	if (mulfprdy = '1') then state := s2670;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2669; end if;
when s2670 => state := s2671; 	--9
	mulfpsclr <= '0';
when s2671 => state := s2672; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2672 => 			--11
	if (mulfprdy = '1') then state := s2673;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2672; end if;
when s2673 => state := s2674; 	--12
	mulfpsclr <= '0';
when s2674 => state := s2675; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2675 => 			--14
	if (addfprdy = '1') then state := s2676;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2675; end if;
when s2676 => state := s2677; 	--15
	addfpsclr <= '0';
when s2677 => state := s2678; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2678 => 			--17
	if (addfprdy = '1') then state := s2679;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2678; end if;
when s2679 => state := s2680; 	--18
	addfpsclr <= '0';
when s2680 => state := s2681; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2681 => 			--20
	if (addfprdy = '1') then state := s2682;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2681; end if;
when s2682 => state := s2683; 	--21
	addfpsclr <= '0';
when s2683 => state := s2684; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (177, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2684 => state := s2685; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (292, 12)); -- offset LSB 244
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s2685 => state := s2686;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (293, 12)); -- offset MSB 245
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2686 => state := s2687; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2687 => 			--4
	if (fixed2floatrdy = '1') then state := s2688;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2687; end if;
when s2688 => state := s2689; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2689 => 			--6
	if (mulfprdy = '1') then state := s2690;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2689; end if;
when s2690 => state := s2691; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2691 => 			--8
	if (mulfprdy = '1') then state := s2692;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2691; end if;
when s2692 => state := s2693; 	--9
	mulfpsclr <= '0';
when s2693 => state := s2694; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2694 => 			--11
	if (mulfprdy = '1') then state := s2695;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2694; end if;
when s2695 => state := s2696; 	--12
	mulfpsclr <= '0';
when s2696 => state := s2697; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2697 => 			--14
	if (addfprdy = '1') then state := s2698;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2697; end if;
when s2698 => state := s2699; 	--15
	addfpsclr <= '0';
when s2699 => state := s2700; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2700 => 			--17
	if (addfprdy = '1') then state := s2701;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2700; end if;
when s2701 => state := s2702; 	--18
	addfpsclr <= '0';
when s2702 => state := s2703; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2703 => 			--20
	if (addfprdy = '1') then state := s2704;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2703; end if;
when s2704 => state := s2705; 	--21
	addfpsclr <= '0';
when s2705 => state := s2706; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (178, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2706 => state := s2707; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (294, 12)); -- offset LSB 246
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s2707 => state := s2708;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (295, 12)); -- offset MSB 247
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2708 => state := s2709; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2709 => 			--4
	if (fixed2floatrdy = '1') then state := s2710;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2709; end if;
when s2710 => state := s2711; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2711 => 			--6
	if (mulfprdy = '1') then state := s2712;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2711; end if;
when s2712 => state := s2713; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2713 => 			--8
	if (mulfprdy = '1') then state := s2714;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2713; end if;
when s2714 => state := s2715; 	--9
	mulfpsclr <= '0';
when s2715 => state := s2716; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2716 => 			--11
	if (mulfprdy = '1') then state := s2717;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2716; end if;
when s2717 => state := s2718; 	--12
	mulfpsclr <= '0';
when s2718 => state := s2719; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2719 => 			--14
	if (addfprdy = '1') then state := s2720;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2719; end if;
when s2720 => state := s2721; 	--15
	addfpsclr <= '0';
when s2721 => state := s2722; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2722 => 			--17
	if (addfprdy = '1') then state := s2723;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2722; end if;
when s2723 => state := s2724; 	--18
	addfpsclr <= '0';
when s2724 => state := s2725; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2725 => 			--20
	if (addfprdy = '1') then state := s2726;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2725; end if;
when s2726 => state := s2727; 	--21
	addfpsclr <= '0';
when s2727 => state := s2728; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (179, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2728 => state := s2729; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (296, 12)); -- offset LSB 248
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s2729 => state := s2730;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (297, 12)); -- offset MSB 249
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2730 => state := s2731; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2731 => 			--4
	if (fixed2floatrdy = '1') then state := s2732;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2731; end if;
when s2732 => state := s2733; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2733 => 			--6
	if (mulfprdy = '1') then state := s2734;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2733; end if;
when s2734 => state := s2735; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2735 => 			--8
	if (mulfprdy = '1') then state := s2736;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2735; end if;
when s2736 => state := s2737; 	--9
	mulfpsclr <= '0';
when s2737 => state := s2738; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2738 => 			--11
	if (mulfprdy = '1') then state := s2739;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2738; end if;
when s2739 => state := s2740; 	--12
	mulfpsclr <= '0';
when s2740 => state := s2741; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2741 => 			--14
	if (addfprdy = '1') then state := s2742;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2741; end if;
when s2742 => state := s2743; 	--15
	addfpsclr <= '0';
when s2743 => state := s2744; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2744 => 			--17
	if (addfprdy = '1') then state := s2745;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2744; end if;
when s2745 => state := s2746; 	--18
	addfpsclr <= '0';
when s2746 => state := s2747; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2747 => 			--20
	if (addfprdy = '1') then state := s2748;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2747; end if;
when s2748 => state := s2749; 	--21
	addfpsclr <= '0';
when s2749 => state := s2750; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (180, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2750 => state := s2751; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (298, 12)); -- offset LSB 250
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s2751 => state := s2752;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (299, 12)); -- offset MSB 251
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2752 => state := s2753; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2753 => 			--4
	if (fixed2floatrdy = '1') then state := s2754;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2753; end if;
when s2754 => state := s2755; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2755 => 			--6
	if (mulfprdy = '1') then state := s2756;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2755; end if;
when s2756 => state := s2757; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2757 => 			--8
	if (mulfprdy = '1') then state := s2758;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2757; end if;
when s2758 => state := s2759; 	--9
	mulfpsclr <= '0';
when s2759 => state := s2760; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2760 => 			--11
	if (mulfprdy = '1') then state := s2761;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2760; end if;
when s2761 => state := s2762; 	--12
	mulfpsclr <= '0';
when s2762 => state := s2763; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2763 => 			--14
	if (addfprdy = '1') then state := s2764;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2763; end if;
when s2764 => state := s2765; 	--15
	addfpsclr <= '0';
when s2765 => state := s2766; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2766 => 			--17
	if (addfprdy = '1') then state := s2767;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2766; end if;
when s2767 => state := s2768; 	--18
	addfpsclr <= '0';
when s2768 => state := s2769; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2769 => 			--20
	if (addfprdy = '1') then state := s2770;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2769; end if;
when s2770 => state := s2771; 	--21
	addfpsclr <= '0';
when s2771 => state := s2772; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (181, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2772 => state := s2773; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (300, 12)); -- offset LSB 252
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s2773 => state := s2774;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (301, 12)); -- offset MSB 253
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2774 => state := s2775; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2775 => 			--4
	if (fixed2floatrdy = '1') then state := s2776;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2775; end if;
when s2776 => state := s2777; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2777 => 			--6
	if (mulfprdy = '1') then state := s2778;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2777; end if;
when s2778 => state := s2779; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2779 => 			--8
	if (mulfprdy = '1') then state := s2780;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2779; end if;
when s2780 => state := s2781; 	--9
	mulfpsclr <= '0';
when s2781 => state := s2782; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2782 => 			--11
	if (mulfprdy = '1') then state := s2783;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2782; end if;
when s2783 => state := s2784; 	--12
	mulfpsclr <= '0';
when s2784 => state := s2785; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2785 => 			--14
	if (addfprdy = '1') then state := s2786;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2785; end if;
when s2786 => state := s2787; 	--15
	addfpsclr <= '0';
when s2787 => state := s2788; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2788 => 			--17
	if (addfprdy = '1') then state := s2789;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2788; end if;
when s2789 => state := s2790; 	--18
	addfpsclr <= '0';
when s2790 => state := s2791; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2791 => 			--20
	if (addfprdy = '1') then state := s2792;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2791; end if;
when s2792 => state := s2793; 	--21
	addfpsclr <= '0';
when s2793 => state := s2794; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (182, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2794 => state := s2795; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (302, 12)); -- offset LSB 254
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s2795 => state := s2796;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (303, 12)); -- offset MSB 255
	addra <= std_logic_vector (to_unsigned (3, 10)); -- OCCrowI 3
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2796 => state := s2797; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2797 => 			--4
	if (fixed2floatrdy = '1') then state := s2798;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2797; end if;
when s2798 => state := s2799; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2799 => 			--6
	if (mulfprdy = '1') then state := s2800;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2799; end if;
when s2800 => state := s2801; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2801 => 			--8
	if (mulfprdy = '1') then state := s2802;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2801; end if;
when s2802 => state := s2803; 	--9
	mulfpsclr <= '0';
when s2803 => state := s2804; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2804 => 			--11
	if (mulfprdy = '1') then state := s2805;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2804; end if;
when s2805 => state := s2806; 	--12
	mulfpsclr <= '0';
when s2806 => state := s2807; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2807 => 			--14
	if (addfprdy = '1') then state := s2808;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2807; end if;
when s2808 => state := s2809; 	--15
	addfpsclr <= '0';
when s2809 => state := s2810; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2810 => 			--17
	if (addfprdy = '1') then state := s2811;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2810; end if;
when s2811 => state := s2812; 	--18
	addfpsclr <= '0';
when s2812 => state := s2813; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2813 => 			--20
	if (addfprdy = '1') then state := s2814;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2813; end if;
when s2814 => state := s2815; 	--21
	addfpsclr <= '0';
when s2815 => state := s2816; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (183, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2816 => state := s2817; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (304, 12)); -- offset LSB 256
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s2817 => state := s2818;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (305, 12)); -- offset MSB 257
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2818 => state := s2819; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2819 => 			--4
	if (fixed2floatrdy = '1') then state := s2820;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2819; end if;
when s2820 => state := s2821; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2821 => 			--6
	if (mulfprdy = '1') then state := s2822;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2821; end if;
when s2822 => state := s2823; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2823 => 			--8
	if (mulfprdy = '1') then state := s2824;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2823; end if;
when s2824 => state := s2825; 	--9
	mulfpsclr <= '0';
when s2825 => state := s2826; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2826 => 			--11
	if (mulfprdy = '1') then state := s2827;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2826; end if;
when s2827 => state := s2828; 	--12
	mulfpsclr <= '0';
when s2828 => state := s2829; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2829 => 			--14
	if (addfprdy = '1') then state := s2830;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2829; end if;
when s2830 => state := s2831; 	--15
	addfpsclr <= '0';
when s2831 => state := s2832; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2832 => 			--17
	if (addfprdy = '1') then state := s2833;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2832; end if;
when s2833 => state := s2834; 	--18
	addfpsclr <= '0';
when s2834 => state := s2835; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2835 => 			--20
	if (addfprdy = '1') then state := s2836;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2835; end if;
when s2836 => state := s2837; 	--21
	addfpsclr <= '0';
when s2837 => state := s2838; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (184, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2838 => state := s2839; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (306, 12)); -- offset LSB 258
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s2839 => state := s2840;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (307, 12)); -- offset MSB 259
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2840 => state := s2841; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2841 => 			--4
	if (fixed2floatrdy = '1') then state := s2842;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2841; end if;
when s2842 => state := s2843; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2843 => 			--6
	if (mulfprdy = '1') then state := s2844;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2843; end if;
when s2844 => state := s2845; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2845 => 			--8
	if (mulfprdy = '1') then state := s2846;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2845; end if;
when s2846 => state := s2847; 	--9
	mulfpsclr <= '0';
when s2847 => state := s2848; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2848 => 			--11
	if (mulfprdy = '1') then state := s2849;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2848; end if;
when s2849 => state := s2850; 	--12
	mulfpsclr <= '0';
when s2850 => state := s2851; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2851 => 			--14
	if (addfprdy = '1') then state := s2852;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2851; end if;
when s2852 => state := s2853; 	--15
	addfpsclr <= '0';
when s2853 => state := s2854; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2854 => 			--17
	if (addfprdy = '1') then state := s2855;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2854; end if;
when s2855 => state := s2856; 	--18
	addfpsclr <= '0';
when s2856 => state := s2857; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2857 => 			--20
	if (addfprdy = '1') then state := s2858;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2857; end if;
when s2858 => state := s2859; 	--21
	addfpsclr <= '0';
when s2859 => state := s2860; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (185, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2860 => state := s2861; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (308, 12)); -- offset LSB 260
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s2861 => state := s2862;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (309, 12)); -- offset MSB 261
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2862 => state := s2863; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2863 => 			--4
	if (fixed2floatrdy = '1') then state := s2864;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2863; end if;
when s2864 => state := s2865; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2865 => 			--6
	if (mulfprdy = '1') then state := s2866;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2865; end if;
when s2866 => state := s2867; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2867 => 			--8
	if (mulfprdy = '1') then state := s2868;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2867; end if;
when s2868 => state := s2869; 	--9
	mulfpsclr <= '0';
when s2869 => state := s2870; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2870 => 			--11
	if (mulfprdy = '1') then state := s2871;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2870; end if;
when s2871 => state := s2872; 	--12
	mulfpsclr <= '0';
when s2872 => state := s2873; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2873 => 			--14
	if (addfprdy = '1') then state := s2874;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2873; end if;
when s2874 => state := s2875; 	--15
	addfpsclr <= '0';
when s2875 => state := s2876; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2876 => 			--17
	if (addfprdy = '1') then state := s2877;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2876; end if;
when s2877 => state := s2878; 	--18
	addfpsclr <= '0';
when s2878 => state := s2879; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2879 => 			--20
	if (addfprdy = '1') then state := s2880;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2879; end if;
when s2880 => state := s2881; 	--21
	addfpsclr <= '0';
when s2881 => state := s2882; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (186, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2882 => state := s2883; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (310, 12)); -- offset LSB 262
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s2883 => state := s2884;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (311, 12)); -- offset MSB 263
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2884 => state := s2885; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2885 => 			--4
	if (fixed2floatrdy = '1') then state := s2886;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2885; end if;
when s2886 => state := s2887; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2887 => 			--6
	if (mulfprdy = '1') then state := s2888;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2887; end if;
when s2888 => state := s2889; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2889 => 			--8
	if (mulfprdy = '1') then state := s2890;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2889; end if;
when s2890 => state := s2891; 	--9
	mulfpsclr <= '0';
when s2891 => state := s2892; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2892 => 			--11
	if (mulfprdy = '1') then state := s2893;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2892; end if;
when s2893 => state := s2894; 	--12
	mulfpsclr <= '0';
when s2894 => state := s2895; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2895 => 			--14
	if (addfprdy = '1') then state := s2896;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2895; end if;
when s2896 => state := s2897; 	--15
	addfpsclr <= '0';
when s2897 => state := s2898; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2898 => 			--17
	if (addfprdy = '1') then state := s2899;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2898; end if;
when s2899 => state := s2900; 	--18
	addfpsclr <= '0';
when s2900 => state := s2901; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2901 => 			--20
	if (addfprdy = '1') then state := s2902;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2901; end if;
when s2902 => state := s2903; 	--21
	addfpsclr <= '0';
when s2903 => state := s2904; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (187, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2904 => state := s2905; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (312, 12)); -- offset LSB 264
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s2905 => state := s2906;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (313, 12)); -- offset MSB 265
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2906 => state := s2907; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2907 => 			--4
	if (fixed2floatrdy = '1') then state := s2908;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2907; end if;
when s2908 => state := s2909; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2909 => 			--6
	if (mulfprdy = '1') then state := s2910;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2909; end if;
when s2910 => state := s2911; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2911 => 			--8
	if (mulfprdy = '1') then state := s2912;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2911; end if;
when s2912 => state := s2913; 	--9
	mulfpsclr <= '0';
when s2913 => state := s2914; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2914 => 			--11
	if (mulfprdy = '1') then state := s2915;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2914; end if;
when s2915 => state := s2916; 	--12
	mulfpsclr <= '0';
when s2916 => state := s2917; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2917 => 			--14
	if (addfprdy = '1') then state := s2918;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2917; end if;
when s2918 => state := s2919; 	--15
	addfpsclr <= '0';
when s2919 => state := s2920; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2920 => 			--17
	if (addfprdy = '1') then state := s2921;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2920; end if;
when s2921 => state := s2922; 	--18
	addfpsclr <= '0';
when s2922 => state := s2923; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2923 => 			--20
	if (addfprdy = '1') then state := s2924;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2923; end if;
when s2924 => state := s2925; 	--21
	addfpsclr <= '0';
when s2925 => state := s2926; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (188, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2926 => state := s2927; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (314, 12)); -- offset LSB 266
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s2927 => state := s2928;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (315, 12)); -- offset MSB 267
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2928 => state := s2929; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2929 => 			--4
	if (fixed2floatrdy = '1') then state := s2930;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2929; end if;
when s2930 => state := s2931; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2931 => 			--6
	if (mulfprdy = '1') then state := s2932;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2931; end if;
when s2932 => state := s2933; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2933 => 			--8
	if (mulfprdy = '1') then state := s2934;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2933; end if;
when s2934 => state := s2935; 	--9
	mulfpsclr <= '0';
when s2935 => state := s2936; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2936 => 			--11
	if (mulfprdy = '1') then state := s2937;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2936; end if;
when s2937 => state := s2938; 	--12
	mulfpsclr <= '0';
when s2938 => state := s2939; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2939 => 			--14
	if (addfprdy = '1') then state := s2940;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2939; end if;
when s2940 => state := s2941; 	--15
	addfpsclr <= '0';
when s2941 => state := s2942; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2942 => 			--17
	if (addfprdy = '1') then state := s2943;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2942; end if;
when s2943 => state := s2944; 	--18
	addfpsclr <= '0';
when s2944 => state := s2945; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2945 => 			--20
	if (addfprdy = '1') then state := s2946;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2945; end if;
when s2946 => state := s2947; 	--21
	addfpsclr <= '0';
when s2947 => state := s2948; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (189, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2948 => state := s2949; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (316, 12)); -- offset LSB 268
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s2949 => state := s2950;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (317, 12)); -- offset MSB 269
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2950 => state := s2951; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2951 => 			--4
	if (fixed2floatrdy = '1') then state := s2952;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2951; end if;
when s2952 => state := s2953; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2953 => 			--6
	if (mulfprdy = '1') then state := s2954;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2953; end if;
when s2954 => state := s2955; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2955 => 			--8
	if (mulfprdy = '1') then state := s2956;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2955; end if;
when s2956 => state := s2957; 	--9
	mulfpsclr <= '0';
when s2957 => state := s2958; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2958 => 			--11
	if (mulfprdy = '1') then state := s2959;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2958; end if;
when s2959 => state := s2960; 	--12
	mulfpsclr <= '0';
when s2960 => state := s2961; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2961 => 			--14
	if (addfprdy = '1') then state := s2962;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2961; end if;
when s2962 => state := s2963; 	--15
	addfpsclr <= '0';
when s2963 => state := s2964; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2964 => 			--17
	if (addfprdy = '1') then state := s2965;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2964; end if;
when s2965 => state := s2966; 	--18
	addfpsclr <= '0';
when s2966 => state := s2967; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2967 => 			--20
	if (addfprdy = '1') then state := s2968;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2967; end if;
when s2968 => state := s2969; 	--21
	addfpsclr <= '0';
when s2969 => state := s2970; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (190, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2970 => state := s2971; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (318, 12)); -- offset LSB 270
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s2971 => state := s2972;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (319, 12)); -- offset MSB 271
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2972 => state := s2973; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2973 => 			--4
	if (fixed2floatrdy = '1') then state := s2974;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2973; end if;
when s2974 => state := s2975; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2975 => 			--6
	if (mulfprdy = '1') then state := s2976;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2975; end if;
when s2976 => state := s2977; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2977 => 			--8
	if (mulfprdy = '1') then state := s2978;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2977; end if;
when s2978 => state := s2979; 	--9
	mulfpsclr <= '0';
when s2979 => state := s2980; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s2980 => 			--11
	if (mulfprdy = '1') then state := s2981;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2980; end if;
when s2981 => state := s2982; 	--12
	mulfpsclr <= '0';
when s2982 => state := s2983; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s2983 => 			--14
	if (addfprdy = '1') then state := s2984;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2983; end if;
when s2984 => state := s2985; 	--15
	addfpsclr <= '0';
when s2985 => state := s2986; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s2986 => 			--17
	if (addfprdy = '1') then state := s2987;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2986; end if;
when s2987 => state := s2988; 	--18
	addfpsclr <= '0';
when s2988 => state := s2989; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s2989 => 			--20
	if (addfprdy = '1') then state := s2990;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s2989; end if;
when s2990 => state := s2991; 	--21
	addfpsclr <= '0';
when s2991 => state := s2992; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (191, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s2992 => state := s2993; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (320, 12)); -- offset LSB 272
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s2993 => state := s2994;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (321, 12)); -- offset MSB 273
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s2994 => state := s2995; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s2995 => 			--4
	if (fixed2floatrdy = '1') then state := s2996;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s2995; end if;
when s2996 => state := s2997; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s2997 => 			--6
	if (mulfprdy = '1') then state := s2998;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2997; end if;
when s2998 => state := s2999; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s2999 => 			--8
	if (mulfprdy = '1') then state := s3000;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s2999; end if;
when s3000 => state := s3001; 	--9
	mulfpsclr <= '0';
when s3001 => state := s3002; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3002 => 			--11
	if (mulfprdy = '1') then state := s3003;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3002; end if;
when s3003 => state := s3004; 	--12
	mulfpsclr <= '0';
when s3004 => state := s3005; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3005 => 			--14
	if (addfprdy = '1') then state := s3006;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3005; end if;
when s3006 => state := s3007; 	--15
	addfpsclr <= '0';
when s3007 => state := s3008; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3008 => 			--17
	if (addfprdy = '1') then state := s3009;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3008; end if;
when s3009 => state := s3010; 	--18
	addfpsclr <= '0';
when s3010 => state := s3011; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3011 => 			--20
	if (addfprdy = '1') then state := s3012;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3011; end if;
when s3012 => state := s3013; 	--21
	addfpsclr <= '0';
when s3013 => state := s3014; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (192, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3014 => state := s3015; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (322, 12)); -- offset LSB 274
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s3015 => state := s3016;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (323, 12)); -- offset MSB 275
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3016 => state := s3017; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3017 => 			--4
	if (fixed2floatrdy = '1') then state := s3018;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3017; end if;
when s3018 => state := s3019; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3019 => 			--6
	if (mulfprdy = '1') then state := s3020;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3019; end if;
when s3020 => state := s3021; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3021 => 			--8
	if (mulfprdy = '1') then state := s3022;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3021; end if;
when s3022 => state := s3023; 	--9
	mulfpsclr <= '0';
when s3023 => state := s3024; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3024 => 			--11
	if (mulfprdy = '1') then state := s3025;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3024; end if;
when s3025 => state := s3026; 	--12
	mulfpsclr <= '0';
when s3026 => state := s3027; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3027 => 			--14
	if (addfprdy = '1') then state := s3028;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3027; end if;
when s3028 => state := s3029; 	--15
	addfpsclr <= '0';
when s3029 => state := s3030; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3030 => 			--17
	if (addfprdy = '1') then state := s3031;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3030; end if;
when s3031 => state := s3032; 	--18
	addfpsclr <= '0';
when s3032 => state := s3033; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3033 => 			--20
	if (addfprdy = '1') then state := s3034;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3033; end if;
when s3034 => state := s3035; 	--21
	addfpsclr <= '0';
when s3035 => state := s3036; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (193, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3036 => state := s3037; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (324, 12)); -- offset LSB 276
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s3037 => state := s3038;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (325, 12)); -- offset MSB 277
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3038 => state := s3039; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3039 => 			--4
	if (fixed2floatrdy = '1') then state := s3040;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3039; end if;
when s3040 => state := s3041; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3041 => 			--6
	if (mulfprdy = '1') then state := s3042;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3041; end if;
when s3042 => state := s3043; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3043 => 			--8
	if (mulfprdy = '1') then state := s3044;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3043; end if;
when s3044 => state := s3045; 	--9
	mulfpsclr <= '0';
when s3045 => state := s3046; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3046 => 			--11
	if (mulfprdy = '1') then state := s3047;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3046; end if;
when s3047 => state := s3048; 	--12
	mulfpsclr <= '0';
when s3048 => state := s3049; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3049 => 			--14
	if (addfprdy = '1') then state := s3050;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3049; end if;
when s3050 => state := s3051; 	--15
	addfpsclr <= '0';
when s3051 => state := s3052; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3052 => 			--17
	if (addfprdy = '1') then state := s3053;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3052; end if;
when s3053 => state := s3054; 	--18
	addfpsclr <= '0';
when s3054 => state := s3055; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3055 => 			--20
	if (addfprdy = '1') then state := s3056;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3055; end if;
when s3056 => state := s3057; 	--21
	addfpsclr <= '0';
when s3057 => state := s3058; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (194, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3058 => state := s3059; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (326, 12)); -- offset LSB 278
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s3059 => state := s3060;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (327, 12)); -- offset MSB 279
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3060 => state := s3061; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3061 => 			--4
	if (fixed2floatrdy = '1') then state := s3062;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3061; end if;
when s3062 => state := s3063; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3063 => 			--6
	if (mulfprdy = '1') then state := s3064;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3063; end if;
when s3064 => state := s3065; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3065 => 			--8
	if (mulfprdy = '1') then state := s3066;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3065; end if;
when s3066 => state := s3067; 	--9
	mulfpsclr <= '0';
when s3067 => state := s3068; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3068 => 			--11
	if (mulfprdy = '1') then state := s3069;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3068; end if;
when s3069 => state := s3070; 	--12
	mulfpsclr <= '0';
when s3070 => state := s3071; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3071 => 			--14
	if (addfprdy = '1') then state := s3072;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3071; end if;
when s3072 => state := s3073; 	--15
	addfpsclr <= '0';
when s3073 => state := s3074; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3074 => 			--17
	if (addfprdy = '1') then state := s3075;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3074; end if;
when s3075 => state := s3076; 	--18
	addfpsclr <= '0';
when s3076 => state := s3077; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3077 => 			--20
	if (addfprdy = '1') then state := s3078;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3077; end if;
when s3078 => state := s3079; 	--21
	addfpsclr <= '0';
when s3079 => state := s3080; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (195, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3080 => state := s3081; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (328, 12)); -- offset LSB 280
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s3081 => state := s3082;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (329, 12)); -- offset MSB 281
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3082 => state := s3083; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3083 => 			--4
	if (fixed2floatrdy = '1') then state := s3084;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3083; end if;
when s3084 => state := s3085; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3085 => 			--6
	if (mulfprdy = '1') then state := s3086;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3085; end if;
when s3086 => state := s3087; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3087 => 			--8
	if (mulfprdy = '1') then state := s3088;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3087; end if;
when s3088 => state := s3089; 	--9
	mulfpsclr <= '0';
when s3089 => state := s3090; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3090 => 			--11
	if (mulfprdy = '1') then state := s3091;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3090; end if;
when s3091 => state := s3092; 	--12
	mulfpsclr <= '0';
when s3092 => state := s3093; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3093 => 			--14
	if (addfprdy = '1') then state := s3094;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3093; end if;
when s3094 => state := s3095; 	--15
	addfpsclr <= '0';
when s3095 => state := s3096; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3096 => 			--17
	if (addfprdy = '1') then state := s3097;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3096; end if;
when s3097 => state := s3098; 	--18
	addfpsclr <= '0';
when s3098 => state := s3099; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3099 => 			--20
	if (addfprdy = '1') then state := s3100;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3099; end if;
when s3100 => state := s3101; 	--21
	addfpsclr <= '0';
when s3101 => state := s3102; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (196, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3102 => state := s3103; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (330, 12)); -- offset LSB 282
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s3103 => state := s3104;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (331, 12)); -- offset MSB 283
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3104 => state := s3105; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3105 => 			--4
	if (fixed2floatrdy = '1') then state := s3106;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3105; end if;
when s3106 => state := s3107; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3107 => 			--6
	if (mulfprdy = '1') then state := s3108;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3107; end if;
when s3108 => state := s3109; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3109 => 			--8
	if (mulfprdy = '1') then state := s3110;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3109; end if;
when s3110 => state := s3111; 	--9
	mulfpsclr <= '0';
when s3111 => state := s3112; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3112 => 			--11
	if (mulfprdy = '1') then state := s3113;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3112; end if;
when s3113 => state := s3114; 	--12
	mulfpsclr <= '0';
when s3114 => state := s3115; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3115 => 			--14
	if (addfprdy = '1') then state := s3116;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3115; end if;
when s3116 => state := s3117; 	--15
	addfpsclr <= '0';
when s3117 => state := s3118; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3118 => 			--17
	if (addfprdy = '1') then state := s3119;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3118; end if;
when s3119 => state := s3120; 	--18
	addfpsclr <= '0';
when s3120 => state := s3121; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3121 => 			--20
	if (addfprdy = '1') then state := s3122;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3121; end if;
when s3122 => state := s3123; 	--21
	addfpsclr <= '0';
when s3123 => state := s3124; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (197, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3124 => state := s3125; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (332, 12)); -- offset LSB 284
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s3125 => state := s3126;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (333, 12)); -- offset MSB 285
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3126 => state := s3127; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3127 => 			--4
	if (fixed2floatrdy = '1') then state := s3128;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3127; end if;
when s3128 => state := s3129; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3129 => 			--6
	if (mulfprdy = '1') then state := s3130;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3129; end if;
when s3130 => state := s3131; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3131 => 			--8
	if (mulfprdy = '1') then state := s3132;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3131; end if;
when s3132 => state := s3133; 	--9
	mulfpsclr <= '0';
when s3133 => state := s3134; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3134 => 			--11
	if (mulfprdy = '1') then state := s3135;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3134; end if;
when s3135 => state := s3136; 	--12
	mulfpsclr <= '0';
when s3136 => state := s3137; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3137 => 			--14
	if (addfprdy = '1') then state := s3138;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3137; end if;
when s3138 => state := s3139; 	--15
	addfpsclr <= '0';
when s3139 => state := s3140; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3140 => 			--17
	if (addfprdy = '1') then state := s3141;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3140; end if;
when s3141 => state := s3142; 	--18
	addfpsclr <= '0';
when s3142 => state := s3143; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3143 => 			--20
	if (addfprdy = '1') then state := s3144;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3143; end if;
when s3144 => state := s3145; 	--21
	addfpsclr <= '0';
when s3145 => state := s3146; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (198, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3146 => state := s3147; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (334, 12)); -- offset LSB 286
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s3147 => state := s3148;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (335, 12)); -- offset MSB 287
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3148 => state := s3149; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3149 => 			--4
	if (fixed2floatrdy = '1') then state := s3150;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3149; end if;
when s3150 => state := s3151; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3151 => 			--6
	if (mulfprdy = '1') then state := s3152;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3151; end if;
when s3152 => state := s3153; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3153 => 			--8
	if (mulfprdy = '1') then state := s3154;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3153; end if;
when s3154 => state := s3155; 	--9
	mulfpsclr <= '0';
when s3155 => state := s3156; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3156 => 			--11
	if (mulfprdy = '1') then state := s3157;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3156; end if;
when s3157 => state := s3158; 	--12
	mulfpsclr <= '0';
when s3158 => state := s3159; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3159 => 			--14
	if (addfprdy = '1') then state := s3160;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3159; end if;
when s3160 => state := s3161; 	--15
	addfpsclr <= '0';
when s3161 => state := s3162; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3162 => 			--17
	if (addfprdy = '1') then state := s3163;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3162; end if;
when s3163 => state := s3164; 	--18
	addfpsclr <= '0';
when s3164 => state := s3165; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3165 => 			--20
	if (addfprdy = '1') then state := s3166;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3165; end if;
when s3166 => state := s3167; 	--21
	addfpsclr <= '0';
when s3167 => state := s3168; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (199, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3168 => state := s3169; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (336, 12)); -- offset LSB 288
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s3169 => state := s3170;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (337, 12)); -- offset MSB 289
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3170 => state := s3171; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3171 => 			--4
	if (fixed2floatrdy = '1') then state := s3172;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3171; end if;
when s3172 => state := s3173; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3173 => 			--6
	if (mulfprdy = '1') then state := s3174;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3173; end if;
when s3174 => state := s3175; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3175 => 			--8
	if (mulfprdy = '1') then state := s3176;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3175; end if;
when s3176 => state := s3177; 	--9
	mulfpsclr <= '0';
when s3177 => state := s3178; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3178 => 			--11
	if (mulfprdy = '1') then state := s3179;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3178; end if;
when s3179 => state := s3180; 	--12
	mulfpsclr <= '0';
when s3180 => state := s3181; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3181 => 			--14
	if (addfprdy = '1') then state := s3182;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3181; end if;
when s3182 => state := s3183; 	--15
	addfpsclr <= '0';
when s3183 => state := s3184; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3184 => 			--17
	if (addfprdy = '1') then state := s3185;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3184; end if;
when s3185 => state := s3186; 	--18
	addfpsclr <= '0';
when s3186 => state := s3187; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3187 => 			--20
	if (addfprdy = '1') then state := s3188;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3187; end if;
when s3188 => state := s3189; 	--21
	addfpsclr <= '0';
when s3189 => state := s3190; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (200, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3190 => state := s3191; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (338, 12)); -- offset LSB 290
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s3191 => state := s3192;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (339, 12)); -- offset MSB 291
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3192 => state := s3193; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3193 => 			--4
	if (fixed2floatrdy = '1') then state := s3194;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3193; end if;
when s3194 => state := s3195; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3195 => 			--6
	if (mulfprdy = '1') then state := s3196;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3195; end if;
when s3196 => state := s3197; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3197 => 			--8
	if (mulfprdy = '1') then state := s3198;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3197; end if;
when s3198 => state := s3199; 	--9
	mulfpsclr <= '0';
when s3199 => state := s3200; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3200 => 			--11
	if (mulfprdy = '1') then state := s3201;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3200; end if;
when s3201 => state := s3202; 	--12
	mulfpsclr <= '0';
when s3202 => state := s3203; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3203 => 			--14
	if (addfprdy = '1') then state := s3204;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3203; end if;
when s3204 => state := s3205; 	--15
	addfpsclr <= '0';
when s3205 => state := s3206; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3206 => 			--17
	if (addfprdy = '1') then state := s3207;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3206; end if;
when s3207 => state := s3208; 	--18
	addfpsclr <= '0';
when s3208 => state := s3209; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3209 => 			--20
	if (addfprdy = '1') then state := s3210;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3209; end if;
when s3210 => state := s3211; 	--21
	addfpsclr <= '0';
when s3211 => state := s3212; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (201, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3212 => state := s3213; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (340, 12)); -- offset LSB 292
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s3213 => state := s3214;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (341, 12)); -- offset MSB 293
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3214 => state := s3215; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3215 => 			--4
	if (fixed2floatrdy = '1') then state := s3216;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3215; end if;
when s3216 => state := s3217; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3217 => 			--6
	if (mulfprdy = '1') then state := s3218;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3217; end if;
when s3218 => state := s3219; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3219 => 			--8
	if (mulfprdy = '1') then state := s3220;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3219; end if;
when s3220 => state := s3221; 	--9
	mulfpsclr <= '0';
when s3221 => state := s3222; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3222 => 			--11
	if (mulfprdy = '1') then state := s3223;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3222; end if;
when s3223 => state := s3224; 	--12
	mulfpsclr <= '0';
when s3224 => state := s3225; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3225 => 			--14
	if (addfprdy = '1') then state := s3226;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3225; end if;
when s3226 => state := s3227; 	--15
	addfpsclr <= '0';
when s3227 => state := s3228; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3228 => 			--17
	if (addfprdy = '1') then state := s3229;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3228; end if;
when s3229 => state := s3230; 	--18
	addfpsclr <= '0';
when s3230 => state := s3231; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3231 => 			--20
	if (addfprdy = '1') then state := s3232;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3231; end if;
when s3232 => state := s3233; 	--21
	addfpsclr <= '0';
when s3233 => state := s3234; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (202, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3234 => state := s3235; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (342, 12)); -- offset LSB 294
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s3235 => state := s3236;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (343, 12)); -- offset MSB 295
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3236 => state := s3237; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3237 => 			--4
	if (fixed2floatrdy = '1') then state := s3238;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3237; end if;
when s3238 => state := s3239; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3239 => 			--6
	if (mulfprdy = '1') then state := s3240;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3239; end if;
when s3240 => state := s3241; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3241 => 			--8
	if (mulfprdy = '1') then state := s3242;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3241; end if;
when s3242 => state := s3243; 	--9
	mulfpsclr <= '0';
when s3243 => state := s3244; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3244 => 			--11
	if (mulfprdy = '1') then state := s3245;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3244; end if;
when s3245 => state := s3246; 	--12
	mulfpsclr <= '0';
when s3246 => state := s3247; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3247 => 			--14
	if (addfprdy = '1') then state := s3248;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3247; end if;
when s3248 => state := s3249; 	--15
	addfpsclr <= '0';
when s3249 => state := s3250; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3250 => 			--17
	if (addfprdy = '1') then state := s3251;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3250; end if;
when s3251 => state := s3252; 	--18
	addfpsclr <= '0';
when s3252 => state := s3253; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3253 => 			--20
	if (addfprdy = '1') then state := s3254;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3253; end if;
when s3254 => state := s3255; 	--21
	addfpsclr <= '0';
when s3255 => state := s3256; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (203, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3256 => state := s3257; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (344, 12)); -- offset LSB 296
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s3257 => state := s3258;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (345, 12)); -- offset MSB 297
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3258 => state := s3259; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3259 => 			--4
	if (fixed2floatrdy = '1') then state := s3260;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3259; end if;
when s3260 => state := s3261; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3261 => 			--6
	if (mulfprdy = '1') then state := s3262;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3261; end if;
when s3262 => state := s3263; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3263 => 			--8
	if (mulfprdy = '1') then state := s3264;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3263; end if;
when s3264 => state := s3265; 	--9
	mulfpsclr <= '0';
when s3265 => state := s3266; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3266 => 			--11
	if (mulfprdy = '1') then state := s3267;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3266; end if;
when s3267 => state := s3268; 	--12
	mulfpsclr <= '0';
when s3268 => state := s3269; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3269 => 			--14
	if (addfprdy = '1') then state := s3270;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3269; end if;
when s3270 => state := s3271; 	--15
	addfpsclr <= '0';
when s3271 => state := s3272; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3272 => 			--17
	if (addfprdy = '1') then state := s3273;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3272; end if;
when s3273 => state := s3274; 	--18
	addfpsclr <= '0';
when s3274 => state := s3275; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3275 => 			--20
	if (addfprdy = '1') then state := s3276;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3275; end if;
when s3276 => state := s3277; 	--21
	addfpsclr <= '0';
when s3277 => state := s3278; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (204, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3278 => state := s3279; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (346, 12)); -- offset LSB 298
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s3279 => state := s3280;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (347, 12)); -- offset MSB 299
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3280 => state := s3281; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3281 => 			--4
	if (fixed2floatrdy = '1') then state := s3282;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3281; end if;
when s3282 => state := s3283; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3283 => 			--6
	if (mulfprdy = '1') then state := s3284;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3283; end if;
when s3284 => state := s3285; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3285 => 			--8
	if (mulfprdy = '1') then state := s3286;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3285; end if;
when s3286 => state := s3287; 	--9
	mulfpsclr <= '0';
when s3287 => state := s3288; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3288 => 			--11
	if (mulfprdy = '1') then state := s3289;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3288; end if;
when s3289 => state := s3290; 	--12
	mulfpsclr <= '0';
when s3290 => state := s3291; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3291 => 			--14
	if (addfprdy = '1') then state := s3292;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3291; end if;
when s3292 => state := s3293; 	--15
	addfpsclr <= '0';
when s3293 => state := s3294; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3294 => 			--17
	if (addfprdy = '1') then state := s3295;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3294; end if;
when s3295 => state := s3296; 	--18
	addfpsclr <= '0';
when s3296 => state := s3297; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3297 => 			--20
	if (addfprdy = '1') then state := s3298;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3297; end if;
when s3298 => state := s3299; 	--21
	addfpsclr <= '0';
when s3299 => state := s3300; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (205, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3300 => state := s3301; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (348, 12)); -- offset LSB 300
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s3301 => state := s3302;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (349, 12)); -- offset MSB 301
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3302 => state := s3303; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3303 => 			--4
	if (fixed2floatrdy = '1') then state := s3304;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3303; end if;
when s3304 => state := s3305; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3305 => 			--6
	if (mulfprdy = '1') then state := s3306;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3305; end if;
when s3306 => state := s3307; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3307 => 			--8
	if (mulfprdy = '1') then state := s3308;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3307; end if;
when s3308 => state := s3309; 	--9
	mulfpsclr <= '0';
when s3309 => state := s3310; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3310 => 			--11
	if (mulfprdy = '1') then state := s3311;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3310; end if;
when s3311 => state := s3312; 	--12
	mulfpsclr <= '0';
when s3312 => state := s3313; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3313 => 			--14
	if (addfprdy = '1') then state := s3314;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3313; end if;
when s3314 => state := s3315; 	--15
	addfpsclr <= '0';
when s3315 => state := s3316; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3316 => 			--17
	if (addfprdy = '1') then state := s3317;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3316; end if;
when s3317 => state := s3318; 	--18
	addfpsclr <= '0';
when s3318 => state := s3319; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3319 => 			--20
	if (addfprdy = '1') then state := s3320;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3319; end if;
when s3320 => state := s3321; 	--21
	addfpsclr <= '0';
when s3321 => state := s3322; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (206, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3322 => state := s3323; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (350, 12)); -- offset LSB 302
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s3323 => state := s3324;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (351, 12)); -- offset MSB 303
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3324 => state := s3325; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3325 => 			--4
	if (fixed2floatrdy = '1') then state := s3326;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3325; end if;
when s3326 => state := s3327; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3327 => 			--6
	if (mulfprdy = '1') then state := s3328;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3327; end if;
when s3328 => state := s3329; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3329 => 			--8
	if (mulfprdy = '1') then state := s3330;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3329; end if;
when s3330 => state := s3331; 	--9
	mulfpsclr <= '0';
when s3331 => state := s3332; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3332 => 			--11
	if (mulfprdy = '1') then state := s3333;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3332; end if;
when s3333 => state := s3334; 	--12
	mulfpsclr <= '0';
when s3334 => state := s3335; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3335 => 			--14
	if (addfprdy = '1') then state := s3336;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3335; end if;
when s3336 => state := s3337; 	--15
	addfpsclr <= '0';
when s3337 => state := s3338; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3338 => 			--17
	if (addfprdy = '1') then state := s3339;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3338; end if;
when s3339 => state := s3340; 	--18
	addfpsclr <= '0';
when s3340 => state := s3341; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3341 => 			--20
	if (addfprdy = '1') then state := s3342;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3341; end if;
when s3342 => state := s3343; 	--21
	addfpsclr <= '0';
when s3343 => state := s3344; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (207, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3344 => state := s3345; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (352, 12)); -- offset LSB 304
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s3345 => state := s3346;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (353, 12)); -- offset MSB 305
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3346 => state := s3347; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3347 => 			--4
	if (fixed2floatrdy = '1') then state := s3348;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3347; end if;
when s3348 => state := s3349; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3349 => 			--6
	if (mulfprdy = '1') then state := s3350;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3349; end if;
when s3350 => state := s3351; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3351 => 			--8
	if (mulfprdy = '1') then state := s3352;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3351; end if;
when s3352 => state := s3353; 	--9
	mulfpsclr <= '0';
when s3353 => state := s3354; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3354 => 			--11
	if (mulfprdy = '1') then state := s3355;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3354; end if;
when s3355 => state := s3356; 	--12
	mulfpsclr <= '0';
when s3356 => state := s3357; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3357 => 			--14
	if (addfprdy = '1') then state := s3358;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3357; end if;
when s3358 => state := s3359; 	--15
	addfpsclr <= '0';
when s3359 => state := s3360; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3360 => 			--17
	if (addfprdy = '1') then state := s3361;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3360; end if;
when s3361 => state := s3362; 	--18
	addfpsclr <= '0';
when s3362 => state := s3363; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3363 => 			--20
	if (addfprdy = '1') then state := s3364;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3363; end if;
when s3364 => state := s3365; 	--21
	addfpsclr <= '0';
when s3365 => state := s3366; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (208, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3366 => state := s3367; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (354, 12)); -- offset LSB 306
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s3367 => state := s3368;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (355, 12)); -- offset MSB 307
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3368 => state := s3369; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3369 => 			--4
	if (fixed2floatrdy = '1') then state := s3370;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3369; end if;
when s3370 => state := s3371; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3371 => 			--6
	if (mulfprdy = '1') then state := s3372;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3371; end if;
when s3372 => state := s3373; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3373 => 			--8
	if (mulfprdy = '1') then state := s3374;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3373; end if;
when s3374 => state := s3375; 	--9
	mulfpsclr <= '0';
when s3375 => state := s3376; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3376 => 			--11
	if (mulfprdy = '1') then state := s3377;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3376; end if;
when s3377 => state := s3378; 	--12
	mulfpsclr <= '0';
when s3378 => state := s3379; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3379 => 			--14
	if (addfprdy = '1') then state := s3380;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3379; end if;
when s3380 => state := s3381; 	--15
	addfpsclr <= '0';
when s3381 => state := s3382; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3382 => 			--17
	if (addfprdy = '1') then state := s3383;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3382; end if;
when s3383 => state := s3384; 	--18
	addfpsclr <= '0';
when s3384 => state := s3385; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3385 => 			--20
	if (addfprdy = '1') then state := s3386;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3385; end if;
when s3386 => state := s3387; 	--21
	addfpsclr <= '0';
when s3387 => state := s3388; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (209, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3388 => state := s3389; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (356, 12)); -- offset LSB 308
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s3389 => state := s3390;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (357, 12)); -- offset MSB 309
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3390 => state := s3391; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3391 => 			--4
	if (fixed2floatrdy = '1') then state := s3392;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3391; end if;
when s3392 => state := s3393; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3393 => 			--6
	if (mulfprdy = '1') then state := s3394;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3393; end if;
when s3394 => state := s3395; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3395 => 			--8
	if (mulfprdy = '1') then state := s3396;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3395; end if;
when s3396 => state := s3397; 	--9
	mulfpsclr <= '0';
when s3397 => state := s3398; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3398 => 			--11
	if (mulfprdy = '1') then state := s3399;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3398; end if;
when s3399 => state := s3400; 	--12
	mulfpsclr <= '0';
when s3400 => state := s3401; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3401 => 			--14
	if (addfprdy = '1') then state := s3402;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3401; end if;
when s3402 => state := s3403; 	--15
	addfpsclr <= '0';
when s3403 => state := s3404; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3404 => 			--17
	if (addfprdy = '1') then state := s3405;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3404; end if;
when s3405 => state := s3406; 	--18
	addfpsclr <= '0';
when s3406 => state := s3407; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3407 => 			--20
	if (addfprdy = '1') then state := s3408;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3407; end if;
when s3408 => state := s3409; 	--21
	addfpsclr <= '0';
when s3409 => state := s3410; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (210, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3410 => state := s3411; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (358, 12)); -- offset LSB 310
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s3411 => state := s3412;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (359, 12)); -- offset MSB 311
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3412 => state := s3413; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3413 => 			--4
	if (fixed2floatrdy = '1') then state := s3414;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3413; end if;
when s3414 => state := s3415; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3415 => 			--6
	if (mulfprdy = '1') then state := s3416;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3415; end if;
when s3416 => state := s3417; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3417 => 			--8
	if (mulfprdy = '1') then state := s3418;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3417; end if;
when s3418 => state := s3419; 	--9
	mulfpsclr <= '0';
when s3419 => state := s3420; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3420 => 			--11
	if (mulfprdy = '1') then state := s3421;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3420; end if;
when s3421 => state := s3422; 	--12
	mulfpsclr <= '0';
when s3422 => state := s3423; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3423 => 			--14
	if (addfprdy = '1') then state := s3424;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3423; end if;
when s3424 => state := s3425; 	--15
	addfpsclr <= '0';
when s3425 => state := s3426; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3426 => 			--17
	if (addfprdy = '1') then state := s3427;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3426; end if;
when s3427 => state := s3428; 	--18
	addfpsclr <= '0';
when s3428 => state := s3429; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3429 => 			--20
	if (addfprdy = '1') then state := s3430;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3429; end if;
when s3430 => state := s3431; 	--21
	addfpsclr <= '0';
when s3431 => state := s3432; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (211, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3432 => state := s3433; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (360, 12)); -- offset LSB 312
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s3433 => state := s3434;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (361, 12)); -- offset MSB 313
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3434 => state := s3435; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3435 => 			--4
	if (fixed2floatrdy = '1') then state := s3436;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3435; end if;
when s3436 => state := s3437; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3437 => 			--6
	if (mulfprdy = '1') then state := s3438;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3437; end if;
when s3438 => state := s3439; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3439 => 			--8
	if (mulfprdy = '1') then state := s3440;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3439; end if;
when s3440 => state := s3441; 	--9
	mulfpsclr <= '0';
when s3441 => state := s3442; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3442 => 			--11
	if (mulfprdy = '1') then state := s3443;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3442; end if;
when s3443 => state := s3444; 	--12
	mulfpsclr <= '0';
when s3444 => state := s3445; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3445 => 			--14
	if (addfprdy = '1') then state := s3446;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3445; end if;
when s3446 => state := s3447; 	--15
	addfpsclr <= '0';
when s3447 => state := s3448; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3448 => 			--17
	if (addfprdy = '1') then state := s3449;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3448; end if;
when s3449 => state := s3450; 	--18
	addfpsclr <= '0';
when s3450 => state := s3451; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3451 => 			--20
	if (addfprdy = '1') then state := s3452;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3451; end if;
when s3452 => state := s3453; 	--21
	addfpsclr <= '0';
when s3453 => state := s3454; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (212, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3454 => state := s3455; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (362, 12)); -- offset LSB 314
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s3455 => state := s3456;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (363, 12)); -- offset MSB 315
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3456 => state := s3457; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3457 => 			--4
	if (fixed2floatrdy = '1') then state := s3458;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3457; end if;
when s3458 => state := s3459; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3459 => 			--6
	if (mulfprdy = '1') then state := s3460;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3459; end if;
when s3460 => state := s3461; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3461 => 			--8
	if (mulfprdy = '1') then state := s3462;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3461; end if;
when s3462 => state := s3463; 	--9
	mulfpsclr <= '0';
when s3463 => state := s3464; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3464 => 			--11
	if (mulfprdy = '1') then state := s3465;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3464; end if;
when s3465 => state := s3466; 	--12
	mulfpsclr <= '0';
when s3466 => state := s3467; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3467 => 			--14
	if (addfprdy = '1') then state := s3468;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3467; end if;
when s3468 => state := s3469; 	--15
	addfpsclr <= '0';
when s3469 => state := s3470; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3470 => 			--17
	if (addfprdy = '1') then state := s3471;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3470; end if;
when s3471 => state := s3472; 	--18
	addfpsclr <= '0';
when s3472 => state := s3473; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3473 => 			--20
	if (addfprdy = '1') then state := s3474;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3473; end if;
when s3474 => state := s3475; 	--21
	addfpsclr <= '0';
when s3475 => state := s3476; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (213, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3476 => state := s3477; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (364, 12)); -- offset LSB 316
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s3477 => state := s3478;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (365, 12)); -- offset MSB 317
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3478 => state := s3479; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3479 => 			--4
	if (fixed2floatrdy = '1') then state := s3480;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3479; end if;
when s3480 => state := s3481; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3481 => 			--6
	if (mulfprdy = '1') then state := s3482;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3481; end if;
when s3482 => state := s3483; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3483 => 			--8
	if (mulfprdy = '1') then state := s3484;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3483; end if;
when s3484 => state := s3485; 	--9
	mulfpsclr <= '0';
when s3485 => state := s3486; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3486 => 			--11
	if (mulfprdy = '1') then state := s3487;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3486; end if;
when s3487 => state := s3488; 	--12
	mulfpsclr <= '0';
when s3488 => state := s3489; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3489 => 			--14
	if (addfprdy = '1') then state := s3490;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3489; end if;
when s3490 => state := s3491; 	--15
	addfpsclr <= '0';
when s3491 => state := s3492; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3492 => 			--17
	if (addfprdy = '1') then state := s3493;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3492; end if;
when s3493 => state := s3494; 	--18
	addfpsclr <= '0';
when s3494 => state := s3495; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3495 => 			--20
	if (addfprdy = '1') then state := s3496;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3495; end if;
when s3496 => state := s3497; 	--21
	addfpsclr <= '0';
when s3497 => state := s3498; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (214, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3498 => state := s3499; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (366, 12)); -- offset LSB 318
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s3499 => state := s3500;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (367, 12)); -- offset MSB 319
	addra <= std_logic_vector (to_unsigned (4, 10)); -- OCCrowI 4
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3500 => state := s3501; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3501 => 			--4
	if (fixed2floatrdy = '1') then state := s3502;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3501; end if;
when s3502 => state := s3503; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3503 => 			--6
	if (mulfprdy = '1') then state := s3504;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3503; end if;
when s3504 => state := s3505; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3505 => 			--8
	if (mulfprdy = '1') then state := s3506;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3505; end if;
when s3506 => state := s3507; 	--9
	mulfpsclr <= '0';
when s3507 => state := s3508; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3508 => 			--11
	if (mulfprdy = '1') then state := s3509;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3508; end if;
when s3509 => state := s3510; 	--12
	mulfpsclr <= '0';
when s3510 => state := s3511; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3511 => 			--14
	if (addfprdy = '1') then state := s3512;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3511; end if;
when s3512 => state := s3513; 	--15
	addfpsclr <= '0';
when s3513 => state := s3514; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3514 => 			--17
	if (addfprdy = '1') then state := s3515;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3514; end if;
when s3515 => state := s3516; 	--18
	addfpsclr <= '0';
when s3516 => state := s3517; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3517 => 			--20
	if (addfprdy = '1') then state := s3518;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3517; end if;
when s3518 => state := s3519; 	--21
	addfpsclr <= '0';
when s3519 => state := s3520; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (215, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3520 => state := s3521; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (368, 12)); -- offset LSB 320
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s3521 => state := s3522;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (369, 12)); -- offset MSB 321
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3522 => state := s3523; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3523 => 			--4
	if (fixed2floatrdy = '1') then state := s3524;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3523; end if;
when s3524 => state := s3525; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3525 => 			--6
	if (mulfprdy = '1') then state := s3526;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3525; end if;
when s3526 => state := s3527; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3527 => 			--8
	if (mulfprdy = '1') then state := s3528;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3527; end if;
when s3528 => state := s3529; 	--9
	mulfpsclr <= '0';
when s3529 => state := s3530; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3530 => 			--11
	if (mulfprdy = '1') then state := s3531;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3530; end if;
when s3531 => state := s3532; 	--12
	mulfpsclr <= '0';
when s3532 => state := s3533; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3533 => 			--14
	if (addfprdy = '1') then state := s3534;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3533; end if;
when s3534 => state := s3535; 	--15
	addfpsclr <= '0';
when s3535 => state := s3536; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3536 => 			--17
	if (addfprdy = '1') then state := s3537;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3536; end if;
when s3537 => state := s3538; 	--18
	addfpsclr <= '0';
when s3538 => state := s3539; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3539 => 			--20
	if (addfprdy = '1') then state := s3540;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3539; end if;
when s3540 => state := s3541; 	--21
	addfpsclr <= '0';
when s3541 => state := s3542; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (216, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3542 => state := s3543; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (370, 12)); -- offset LSB 322
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s3543 => state := s3544;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (371, 12)); -- offset MSB 323
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3544 => state := s3545; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3545 => 			--4
	if (fixed2floatrdy = '1') then state := s3546;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3545; end if;
when s3546 => state := s3547; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3547 => 			--6
	if (mulfprdy = '1') then state := s3548;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3547; end if;
when s3548 => state := s3549; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3549 => 			--8
	if (mulfprdy = '1') then state := s3550;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3549; end if;
when s3550 => state := s3551; 	--9
	mulfpsclr <= '0';
when s3551 => state := s3552; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3552 => 			--11
	if (mulfprdy = '1') then state := s3553;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3552; end if;
when s3553 => state := s3554; 	--12
	mulfpsclr <= '0';
when s3554 => state := s3555; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3555 => 			--14
	if (addfprdy = '1') then state := s3556;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3555; end if;
when s3556 => state := s3557; 	--15
	addfpsclr <= '0';
when s3557 => state := s3558; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3558 => 			--17
	if (addfprdy = '1') then state := s3559;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3558; end if;
when s3559 => state := s3560; 	--18
	addfpsclr <= '0';
when s3560 => state := s3561; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3561 => 			--20
	if (addfprdy = '1') then state := s3562;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3561; end if;
when s3562 => state := s3563; 	--21
	addfpsclr <= '0';
when s3563 => state := s3564; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (217, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3564 => state := s3565; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (372, 12)); -- offset LSB 324
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s3565 => state := s3566;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (373, 12)); -- offset MSB 325
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3566 => state := s3567; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3567 => 			--4
	if (fixed2floatrdy = '1') then state := s3568;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3567; end if;
when s3568 => state := s3569; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3569 => 			--6
	if (mulfprdy = '1') then state := s3570;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3569; end if;
when s3570 => state := s3571; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3571 => 			--8
	if (mulfprdy = '1') then state := s3572;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3571; end if;
when s3572 => state := s3573; 	--9
	mulfpsclr <= '0';
when s3573 => state := s3574; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3574 => 			--11
	if (mulfprdy = '1') then state := s3575;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3574; end if;
when s3575 => state := s3576; 	--12
	mulfpsclr <= '0';
when s3576 => state := s3577; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3577 => 			--14
	if (addfprdy = '1') then state := s3578;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3577; end if;
when s3578 => state := s3579; 	--15
	addfpsclr <= '0';
when s3579 => state := s3580; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3580 => 			--17
	if (addfprdy = '1') then state := s3581;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3580; end if;
when s3581 => state := s3582; 	--18
	addfpsclr <= '0';
when s3582 => state := s3583; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3583 => 			--20
	if (addfprdy = '1') then state := s3584;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3583; end if;
when s3584 => state := s3585; 	--21
	addfpsclr <= '0';
when s3585 => state := s3586; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (218, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3586 => state := s3587; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (374, 12)); -- offset LSB 326
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s3587 => state := s3588;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (375, 12)); -- offset MSB 327
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3588 => state := s3589; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3589 => 			--4
	if (fixed2floatrdy = '1') then state := s3590;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3589; end if;
when s3590 => state := s3591; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3591 => 			--6
	if (mulfprdy = '1') then state := s3592;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3591; end if;
when s3592 => state := s3593; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3593 => 			--8
	if (mulfprdy = '1') then state := s3594;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3593; end if;
when s3594 => state := s3595; 	--9
	mulfpsclr <= '0';
when s3595 => state := s3596; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3596 => 			--11
	if (mulfprdy = '1') then state := s3597;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3596; end if;
when s3597 => state := s3598; 	--12
	mulfpsclr <= '0';
when s3598 => state := s3599; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3599 => 			--14
	if (addfprdy = '1') then state := s3600;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3599; end if;
when s3600 => state := s3601; 	--15
	addfpsclr <= '0';
when s3601 => state := s3602; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3602 => 			--17
	if (addfprdy = '1') then state := s3603;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3602; end if;
when s3603 => state := s3604; 	--18
	addfpsclr <= '0';
when s3604 => state := s3605; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3605 => 			--20
	if (addfprdy = '1') then state := s3606;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3605; end if;
when s3606 => state := s3607; 	--21
	addfpsclr <= '0';
when s3607 => state := s3608; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (219, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3608 => state := s3609; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (376, 12)); -- offset LSB 328
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s3609 => state := s3610;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (377, 12)); -- offset MSB 329
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3610 => state := s3611; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3611 => 			--4
	if (fixed2floatrdy = '1') then state := s3612;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3611; end if;
when s3612 => state := s3613; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3613 => 			--6
	if (mulfprdy = '1') then state := s3614;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3613; end if;
when s3614 => state := s3615; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3615 => 			--8
	if (mulfprdy = '1') then state := s3616;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3615; end if;
when s3616 => state := s3617; 	--9
	mulfpsclr <= '0';
when s3617 => state := s3618; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3618 => 			--11
	if (mulfprdy = '1') then state := s3619;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3618; end if;
when s3619 => state := s3620; 	--12
	mulfpsclr <= '0';
when s3620 => state := s3621; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3621 => 			--14
	if (addfprdy = '1') then state := s3622;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3621; end if;
when s3622 => state := s3623; 	--15
	addfpsclr <= '0';
when s3623 => state := s3624; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3624 => 			--17
	if (addfprdy = '1') then state := s3625;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3624; end if;
when s3625 => state := s3626; 	--18
	addfpsclr <= '0';
when s3626 => state := s3627; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3627 => 			--20
	if (addfprdy = '1') then state := s3628;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3627; end if;
when s3628 => state := s3629; 	--21
	addfpsclr <= '0';
when s3629 => state := s3630; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (220, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3630 => state := s3631; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (378, 12)); -- offset LSB 330
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s3631 => state := s3632;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (379, 12)); -- offset MSB 331
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3632 => state := s3633; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3633 => 			--4
	if (fixed2floatrdy = '1') then state := s3634;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3633; end if;
when s3634 => state := s3635; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3635 => 			--6
	if (mulfprdy = '1') then state := s3636;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3635; end if;
when s3636 => state := s3637; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3637 => 			--8
	if (mulfprdy = '1') then state := s3638;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3637; end if;
when s3638 => state := s3639; 	--9
	mulfpsclr <= '0';
when s3639 => state := s3640; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3640 => 			--11
	if (mulfprdy = '1') then state := s3641;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3640; end if;
when s3641 => state := s3642; 	--12
	mulfpsclr <= '0';
when s3642 => state := s3643; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3643 => 			--14
	if (addfprdy = '1') then state := s3644;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3643; end if;
when s3644 => state := s3645; 	--15
	addfpsclr <= '0';
when s3645 => state := s3646; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3646 => 			--17
	if (addfprdy = '1') then state := s3647;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3646; end if;
when s3647 => state := s3648; 	--18
	addfpsclr <= '0';
when s3648 => state := s3649; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3649 => 			--20
	if (addfprdy = '1') then state := s3650;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3649; end if;
when s3650 => state := s3651; 	--21
	addfpsclr <= '0';
when s3651 => state := s3652; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (221, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3652 => state := s3653; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (380, 12)); -- offset LSB 332
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s3653 => state := s3654;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (381, 12)); -- offset MSB 333
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3654 => state := s3655; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3655 => 			--4
	if (fixed2floatrdy = '1') then state := s3656;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3655; end if;
when s3656 => state := s3657; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3657 => 			--6
	if (mulfprdy = '1') then state := s3658;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3657; end if;
when s3658 => state := s3659; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3659 => 			--8
	if (mulfprdy = '1') then state := s3660;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3659; end if;
when s3660 => state := s3661; 	--9
	mulfpsclr <= '0';
when s3661 => state := s3662; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3662 => 			--11
	if (mulfprdy = '1') then state := s3663;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3662; end if;
when s3663 => state := s3664; 	--12
	mulfpsclr <= '0';
when s3664 => state := s3665; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3665 => 			--14
	if (addfprdy = '1') then state := s3666;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3665; end if;
when s3666 => state := s3667; 	--15
	addfpsclr <= '0';
when s3667 => state := s3668; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3668 => 			--17
	if (addfprdy = '1') then state := s3669;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3668; end if;
when s3669 => state := s3670; 	--18
	addfpsclr <= '0';
when s3670 => state := s3671; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3671 => 			--20
	if (addfprdy = '1') then state := s3672;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3671; end if;
when s3672 => state := s3673; 	--21
	addfpsclr <= '0';
when s3673 => state := s3674; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (222, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3674 => state := s3675; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (382, 12)); -- offset LSB 334
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s3675 => state := s3676;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (383, 12)); -- offset MSB 335
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3676 => state := s3677; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3677 => 			--4
	if (fixed2floatrdy = '1') then state := s3678;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3677; end if;
when s3678 => state := s3679; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3679 => 			--6
	if (mulfprdy = '1') then state := s3680;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3679; end if;
when s3680 => state := s3681; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3681 => 			--8
	if (mulfprdy = '1') then state := s3682;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3681; end if;
when s3682 => state := s3683; 	--9
	mulfpsclr <= '0';
when s3683 => state := s3684; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3684 => 			--11
	if (mulfprdy = '1') then state := s3685;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3684; end if;
when s3685 => state := s3686; 	--12
	mulfpsclr <= '0';
when s3686 => state := s3687; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3687 => 			--14
	if (addfprdy = '1') then state := s3688;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3687; end if;
when s3688 => state := s3689; 	--15
	addfpsclr <= '0';
when s3689 => state := s3690; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3690 => 			--17
	if (addfprdy = '1') then state := s3691;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3690; end if;
when s3691 => state := s3692; 	--18
	addfpsclr <= '0';
when s3692 => state := s3693; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3693 => 			--20
	if (addfprdy = '1') then state := s3694;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3693; end if;
when s3694 => state := s3695; 	--21
	addfpsclr <= '0';
when s3695 => state := s3696; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (223, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3696 => state := s3697; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (384, 12)); -- offset LSB 336
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s3697 => state := s3698;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (385, 12)); -- offset MSB 337
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3698 => state := s3699; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3699 => 			--4
	if (fixed2floatrdy = '1') then state := s3700;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3699; end if;
when s3700 => state := s3701; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3701 => 			--6
	if (mulfprdy = '1') then state := s3702;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3701; end if;
when s3702 => state := s3703; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3703 => 			--8
	if (mulfprdy = '1') then state := s3704;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3703; end if;
when s3704 => state := s3705; 	--9
	mulfpsclr <= '0';
when s3705 => state := s3706; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3706 => 			--11
	if (mulfprdy = '1') then state := s3707;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3706; end if;
when s3707 => state := s3708; 	--12
	mulfpsclr <= '0';
when s3708 => state := s3709; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3709 => 			--14
	if (addfprdy = '1') then state := s3710;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3709; end if;
when s3710 => state := s3711; 	--15
	addfpsclr <= '0';
when s3711 => state := s3712; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3712 => 			--17
	if (addfprdy = '1') then state := s3713;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3712; end if;
when s3713 => state := s3714; 	--18
	addfpsclr <= '0';
when s3714 => state := s3715; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3715 => 			--20
	if (addfprdy = '1') then state := s3716;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3715; end if;
when s3716 => state := s3717; 	--21
	addfpsclr <= '0';
when s3717 => state := s3718; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (224, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3718 => state := s3719; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (386, 12)); -- offset LSB 338
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s3719 => state := s3720;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (387, 12)); -- offset MSB 339
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3720 => state := s3721; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3721 => 			--4
	if (fixed2floatrdy = '1') then state := s3722;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3721; end if;
when s3722 => state := s3723; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3723 => 			--6
	if (mulfprdy = '1') then state := s3724;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3723; end if;
when s3724 => state := s3725; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3725 => 			--8
	if (mulfprdy = '1') then state := s3726;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3725; end if;
when s3726 => state := s3727; 	--9
	mulfpsclr <= '0';
when s3727 => state := s3728; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3728 => 			--11
	if (mulfprdy = '1') then state := s3729;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3728; end if;
when s3729 => state := s3730; 	--12
	mulfpsclr <= '0';
when s3730 => state := s3731; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3731 => 			--14
	if (addfprdy = '1') then state := s3732;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3731; end if;
when s3732 => state := s3733; 	--15
	addfpsclr <= '0';
when s3733 => state := s3734; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3734 => 			--17
	if (addfprdy = '1') then state := s3735;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3734; end if;
when s3735 => state := s3736; 	--18
	addfpsclr <= '0';
when s3736 => state := s3737; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3737 => 			--20
	if (addfprdy = '1') then state := s3738;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3737; end if;
when s3738 => state := s3739; 	--21
	addfpsclr <= '0';
when s3739 => state := s3740; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (225, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3740 => state := s3741; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (388, 12)); -- offset LSB 340
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s3741 => state := s3742;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (389, 12)); -- offset MSB 341
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3742 => state := s3743; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3743 => 			--4
	if (fixed2floatrdy = '1') then state := s3744;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3743; end if;
when s3744 => state := s3745; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3745 => 			--6
	if (mulfprdy = '1') then state := s3746;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3745; end if;
when s3746 => state := s3747; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3747 => 			--8
	if (mulfprdy = '1') then state := s3748;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3747; end if;
when s3748 => state := s3749; 	--9
	mulfpsclr <= '0';
when s3749 => state := s3750; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3750 => 			--11
	if (mulfprdy = '1') then state := s3751;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3750; end if;
when s3751 => state := s3752; 	--12
	mulfpsclr <= '0';
when s3752 => state := s3753; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3753 => 			--14
	if (addfprdy = '1') then state := s3754;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3753; end if;
when s3754 => state := s3755; 	--15
	addfpsclr <= '0';
when s3755 => state := s3756; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3756 => 			--17
	if (addfprdy = '1') then state := s3757;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3756; end if;
when s3757 => state := s3758; 	--18
	addfpsclr <= '0';
when s3758 => state := s3759; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3759 => 			--20
	if (addfprdy = '1') then state := s3760;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3759; end if;
when s3760 => state := s3761; 	--21
	addfpsclr <= '0';
when s3761 => state := s3762; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (226, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3762 => state := s3763; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (390, 12)); -- offset LSB 342
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s3763 => state := s3764;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (391, 12)); -- offset MSB 343
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3764 => state := s3765; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3765 => 			--4
	if (fixed2floatrdy = '1') then state := s3766;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3765; end if;
when s3766 => state := s3767; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3767 => 			--6
	if (mulfprdy = '1') then state := s3768;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3767; end if;
when s3768 => state := s3769; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3769 => 			--8
	if (mulfprdy = '1') then state := s3770;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3769; end if;
when s3770 => state := s3771; 	--9
	mulfpsclr <= '0';
when s3771 => state := s3772; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3772 => 			--11
	if (mulfprdy = '1') then state := s3773;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3772; end if;
when s3773 => state := s3774; 	--12
	mulfpsclr <= '0';
when s3774 => state := s3775; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3775 => 			--14
	if (addfprdy = '1') then state := s3776;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3775; end if;
when s3776 => state := s3777; 	--15
	addfpsclr <= '0';
when s3777 => state := s3778; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3778 => 			--17
	if (addfprdy = '1') then state := s3779;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3778; end if;
when s3779 => state := s3780; 	--18
	addfpsclr <= '0';
when s3780 => state := s3781; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3781 => 			--20
	if (addfprdy = '1') then state := s3782;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3781; end if;
when s3782 => state := s3783; 	--21
	addfpsclr <= '0';
when s3783 => state := s3784; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (227, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3784 => state := s3785; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (392, 12)); -- offset LSB 344
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s3785 => state := s3786;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (393, 12)); -- offset MSB 345
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3786 => state := s3787; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3787 => 			--4
	if (fixed2floatrdy = '1') then state := s3788;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3787; end if;
when s3788 => state := s3789; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3789 => 			--6
	if (mulfprdy = '1') then state := s3790;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3789; end if;
when s3790 => state := s3791; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3791 => 			--8
	if (mulfprdy = '1') then state := s3792;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3791; end if;
when s3792 => state := s3793; 	--9
	mulfpsclr <= '0';
when s3793 => state := s3794; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3794 => 			--11
	if (mulfprdy = '1') then state := s3795;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3794; end if;
when s3795 => state := s3796; 	--12
	mulfpsclr <= '0';
when s3796 => state := s3797; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3797 => 			--14
	if (addfprdy = '1') then state := s3798;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3797; end if;
when s3798 => state := s3799; 	--15
	addfpsclr <= '0';
when s3799 => state := s3800; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3800 => 			--17
	if (addfprdy = '1') then state := s3801;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3800; end if;
when s3801 => state := s3802; 	--18
	addfpsclr <= '0';
when s3802 => state := s3803; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3803 => 			--20
	if (addfprdy = '1') then state := s3804;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3803; end if;
when s3804 => state := s3805; 	--21
	addfpsclr <= '0';
when s3805 => state := s3806; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (228, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3806 => state := s3807; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (394, 12)); -- offset LSB 346
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s3807 => state := s3808;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (395, 12)); -- offset MSB 347
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3808 => state := s3809; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3809 => 			--4
	if (fixed2floatrdy = '1') then state := s3810;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3809; end if;
when s3810 => state := s3811; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3811 => 			--6
	if (mulfprdy = '1') then state := s3812;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3811; end if;
when s3812 => state := s3813; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3813 => 			--8
	if (mulfprdy = '1') then state := s3814;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3813; end if;
when s3814 => state := s3815; 	--9
	mulfpsclr <= '0';
when s3815 => state := s3816; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3816 => 			--11
	if (mulfprdy = '1') then state := s3817;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3816; end if;
when s3817 => state := s3818; 	--12
	mulfpsclr <= '0';
when s3818 => state := s3819; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3819 => 			--14
	if (addfprdy = '1') then state := s3820;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3819; end if;
when s3820 => state := s3821; 	--15
	addfpsclr <= '0';
when s3821 => state := s3822; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3822 => 			--17
	if (addfprdy = '1') then state := s3823;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3822; end if;
when s3823 => state := s3824; 	--18
	addfpsclr <= '0';
when s3824 => state := s3825; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3825 => 			--20
	if (addfprdy = '1') then state := s3826;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3825; end if;
when s3826 => state := s3827; 	--21
	addfpsclr <= '0';
when s3827 => state := s3828; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (229, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3828 => state := s3829; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (396, 12)); -- offset LSB 348
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s3829 => state := s3830;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (397, 12)); -- offset MSB 349
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3830 => state := s3831; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3831 => 			--4
	if (fixed2floatrdy = '1') then state := s3832;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3831; end if;
when s3832 => state := s3833; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3833 => 			--6
	if (mulfprdy = '1') then state := s3834;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3833; end if;
when s3834 => state := s3835; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3835 => 			--8
	if (mulfprdy = '1') then state := s3836;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3835; end if;
when s3836 => state := s3837; 	--9
	mulfpsclr <= '0';
when s3837 => state := s3838; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3838 => 			--11
	if (mulfprdy = '1') then state := s3839;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3838; end if;
when s3839 => state := s3840; 	--12
	mulfpsclr <= '0';
when s3840 => state := s3841; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3841 => 			--14
	if (addfprdy = '1') then state := s3842;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3841; end if;
when s3842 => state := s3843; 	--15
	addfpsclr <= '0';
when s3843 => state := s3844; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3844 => 			--17
	if (addfprdy = '1') then state := s3845;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3844; end if;
when s3845 => state := s3846; 	--18
	addfpsclr <= '0';
when s3846 => state := s3847; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3847 => 			--20
	if (addfprdy = '1') then state := s3848;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3847; end if;
when s3848 => state := s3849; 	--21
	addfpsclr <= '0';
when s3849 => state := s3850; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (230, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3850 => state := s3851; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (398, 12)); -- offset LSB 350
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s3851 => state := s3852;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (399, 12)); -- offset MSB 351
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3852 => state := s3853; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3853 => 			--4
	if (fixed2floatrdy = '1') then state := s3854;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3853; end if;
when s3854 => state := s3855; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3855 => 			--6
	if (mulfprdy = '1') then state := s3856;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3855; end if;
when s3856 => state := s3857; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3857 => 			--8
	if (mulfprdy = '1') then state := s3858;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3857; end if;
when s3858 => state := s3859; 	--9
	mulfpsclr <= '0';
when s3859 => state := s3860; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3860 => 			--11
	if (mulfprdy = '1') then state := s3861;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3860; end if;
when s3861 => state := s3862; 	--12
	mulfpsclr <= '0';
when s3862 => state := s3863; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3863 => 			--14
	if (addfprdy = '1') then state := s3864;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3863; end if;
when s3864 => state := s3865; 	--15
	addfpsclr <= '0';
when s3865 => state := s3866; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3866 => 			--17
	if (addfprdy = '1') then state := s3867;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3866; end if;
when s3867 => state := s3868; 	--18
	addfpsclr <= '0';
when s3868 => state := s3869; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3869 => 			--20
	if (addfprdy = '1') then state := s3870;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3869; end if;
when s3870 => state := s3871; 	--21
	addfpsclr <= '0';
when s3871 => state := s3872; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (231, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3872 => state := s3873; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (400, 12)); -- offset LSB 352
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s3873 => state := s3874;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (401, 12)); -- offset MSB 353
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3874 => state := s3875; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3875 => 			--4
	if (fixed2floatrdy = '1') then state := s3876;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3875; end if;
when s3876 => state := s3877; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3877 => 			--6
	if (mulfprdy = '1') then state := s3878;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3877; end if;
when s3878 => state := s3879; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3879 => 			--8
	if (mulfprdy = '1') then state := s3880;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3879; end if;
when s3880 => state := s3881; 	--9
	mulfpsclr <= '0';
when s3881 => state := s3882; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3882 => 			--11
	if (mulfprdy = '1') then state := s3883;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3882; end if;
when s3883 => state := s3884; 	--12
	mulfpsclr <= '0';
when s3884 => state := s3885; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3885 => 			--14
	if (addfprdy = '1') then state := s3886;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3885; end if;
when s3886 => state := s3887; 	--15
	addfpsclr <= '0';
when s3887 => state := s3888; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3888 => 			--17
	if (addfprdy = '1') then state := s3889;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3888; end if;
when s3889 => state := s3890; 	--18
	addfpsclr <= '0';
when s3890 => state := s3891; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3891 => 			--20
	if (addfprdy = '1') then state := s3892;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3891; end if;
when s3892 => state := s3893; 	--21
	addfpsclr <= '0';
when s3893 => state := s3894; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (232, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3894 => state := s3895; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (402, 12)); -- offset LSB 354
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s3895 => state := s3896;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (403, 12)); -- offset MSB 355
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3896 => state := s3897; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3897 => 			--4
	if (fixed2floatrdy = '1') then state := s3898;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3897; end if;
when s3898 => state := s3899; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3899 => 			--6
	if (mulfprdy = '1') then state := s3900;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3899; end if;
when s3900 => state := s3901; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3901 => 			--8
	if (mulfprdy = '1') then state := s3902;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3901; end if;
when s3902 => state := s3903; 	--9
	mulfpsclr <= '0';
when s3903 => state := s3904; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3904 => 			--11
	if (mulfprdy = '1') then state := s3905;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3904; end if;
when s3905 => state := s3906; 	--12
	mulfpsclr <= '0';
when s3906 => state := s3907; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3907 => 			--14
	if (addfprdy = '1') then state := s3908;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3907; end if;
when s3908 => state := s3909; 	--15
	addfpsclr <= '0';
when s3909 => state := s3910; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3910 => 			--17
	if (addfprdy = '1') then state := s3911;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3910; end if;
when s3911 => state := s3912; 	--18
	addfpsclr <= '0';
when s3912 => state := s3913; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3913 => 			--20
	if (addfprdy = '1') then state := s3914;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3913; end if;
when s3914 => state := s3915; 	--21
	addfpsclr <= '0';
when s3915 => state := s3916; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (233, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3916 => state := s3917; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (404, 12)); -- offset LSB 356
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s3917 => state := s3918;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (405, 12)); -- offset MSB 357
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3918 => state := s3919; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3919 => 			--4
	if (fixed2floatrdy = '1') then state := s3920;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3919; end if;
when s3920 => state := s3921; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3921 => 			--6
	if (mulfprdy = '1') then state := s3922;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3921; end if;
when s3922 => state := s3923; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3923 => 			--8
	if (mulfprdy = '1') then state := s3924;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3923; end if;
when s3924 => state := s3925; 	--9
	mulfpsclr <= '0';
when s3925 => state := s3926; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3926 => 			--11
	if (mulfprdy = '1') then state := s3927;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3926; end if;
when s3927 => state := s3928; 	--12
	mulfpsclr <= '0';
when s3928 => state := s3929; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3929 => 			--14
	if (addfprdy = '1') then state := s3930;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3929; end if;
when s3930 => state := s3931; 	--15
	addfpsclr <= '0';
when s3931 => state := s3932; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3932 => 			--17
	if (addfprdy = '1') then state := s3933;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3932; end if;
when s3933 => state := s3934; 	--18
	addfpsclr <= '0';
when s3934 => state := s3935; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3935 => 			--20
	if (addfprdy = '1') then state := s3936;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3935; end if;
when s3936 => state := s3937; 	--21
	addfpsclr <= '0';
when s3937 => state := s3938; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (234, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3938 => state := s3939; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (406, 12)); -- offset LSB 358
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s3939 => state := s3940;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (407, 12)); -- offset MSB 359
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3940 => state := s3941; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3941 => 			--4
	if (fixed2floatrdy = '1') then state := s3942;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3941; end if;
when s3942 => state := s3943; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3943 => 			--6
	if (mulfprdy = '1') then state := s3944;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3943; end if;
when s3944 => state := s3945; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3945 => 			--8
	if (mulfprdy = '1') then state := s3946;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3945; end if;
when s3946 => state := s3947; 	--9
	mulfpsclr <= '0';
when s3947 => state := s3948; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3948 => 			--11
	if (mulfprdy = '1') then state := s3949;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3948; end if;
when s3949 => state := s3950; 	--12
	mulfpsclr <= '0';
when s3950 => state := s3951; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3951 => 			--14
	if (addfprdy = '1') then state := s3952;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3951; end if;
when s3952 => state := s3953; 	--15
	addfpsclr <= '0';
when s3953 => state := s3954; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3954 => 			--17
	if (addfprdy = '1') then state := s3955;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3954; end if;
when s3955 => state := s3956; 	--18
	addfpsclr <= '0';
when s3956 => state := s3957; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3957 => 			--20
	if (addfprdy = '1') then state := s3958;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3957; end if;
when s3958 => state := s3959; 	--21
	addfpsclr <= '0';
when s3959 => state := s3960; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (235, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3960 => state := s3961; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (408, 12)); -- offset LSB 360
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s3961 => state := s3962;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (409, 12)); -- offset MSB 361
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3962 => state := s3963; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3963 => 			--4
	if (fixed2floatrdy = '1') then state := s3964;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3963; end if;
when s3964 => state := s3965; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3965 => 			--6
	if (mulfprdy = '1') then state := s3966;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3965; end if;
when s3966 => state := s3967; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3967 => 			--8
	if (mulfprdy = '1') then state := s3968;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3967; end if;
when s3968 => state := s3969; 	--9
	mulfpsclr <= '0';
when s3969 => state := s3970; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3970 => 			--11
	if (mulfprdy = '1') then state := s3971;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3970; end if;
when s3971 => state := s3972; 	--12
	mulfpsclr <= '0';
when s3972 => state := s3973; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3973 => 			--14
	if (addfprdy = '1') then state := s3974;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3973; end if;
when s3974 => state := s3975; 	--15
	addfpsclr <= '0';
when s3975 => state := s3976; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3976 => 			--17
	if (addfprdy = '1') then state := s3977;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3976; end if;
when s3977 => state := s3978; 	--18
	addfpsclr <= '0';
when s3978 => state := s3979; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s3979 => 			--20
	if (addfprdy = '1') then state := s3980;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3979; end if;
when s3980 => state := s3981; 	--21
	addfpsclr <= '0';
when s3981 => state := s3982; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (236, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s3982 => state := s3983; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (410, 12)); -- offset LSB 362
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s3983 => state := s3984;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (411, 12)); -- offset MSB 363
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s3984 => state := s3985; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s3985 => 			--4
	if (fixed2floatrdy = '1') then state := s3986;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s3985; end if;
when s3986 => state := s3987; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s3987 => 			--6
	if (mulfprdy = '1') then state := s3988;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3987; end if;
when s3988 => state := s3989; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s3989 => 			--8
	if (mulfprdy = '1') then state := s3990;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3989; end if;
when s3990 => state := s3991; 	--9
	mulfpsclr <= '0';
when s3991 => state := s3992; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s3992 => 			--11
	if (mulfprdy = '1') then state := s3993;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s3992; end if;
when s3993 => state := s3994; 	--12
	mulfpsclr <= '0';
when s3994 => state := s3995; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s3995 => 			--14
	if (addfprdy = '1') then state := s3996;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3995; end if;
when s3996 => state := s3997; 	--15
	addfpsclr <= '0';
when s3997 => state := s3998; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s3998 => 			--17
	if (addfprdy = '1') then state := s3999;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s3998; end if;
when s3999 => state := s4000; 	--18
	addfpsclr <= '0';
when s4000 => state := s4001; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4001 => 			--20
	if (addfprdy = '1') then state := s4002;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4001; end if;
when s4002 => state := s4003; 	--21
	addfpsclr <= '0';
when s4003 => state := s4004; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (237, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4004 => state := s4005; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (412, 12)); -- offset LSB 364
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s4005 => state := s4006;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (413, 12)); -- offset MSB 365
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4006 => state := s4007; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4007 => 			--4
	if (fixed2floatrdy = '1') then state := s4008;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4007; end if;
when s4008 => state := s4009; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4009 => 			--6
	if (mulfprdy = '1') then state := s4010;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4009; end if;
when s4010 => state := s4011; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4011 => 			--8
	if (mulfprdy = '1') then state := s4012;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4011; end if;
when s4012 => state := s4013; 	--9
	mulfpsclr <= '0';
when s4013 => state := s4014; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4014 => 			--11
	if (mulfprdy = '1') then state := s4015;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4014; end if;
when s4015 => state := s4016; 	--12
	mulfpsclr <= '0';
when s4016 => state := s4017; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4017 => 			--14
	if (addfprdy = '1') then state := s4018;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4017; end if;
when s4018 => state := s4019; 	--15
	addfpsclr <= '0';
when s4019 => state := s4020; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4020 => 			--17
	if (addfprdy = '1') then state := s4021;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4020; end if;
when s4021 => state := s4022; 	--18
	addfpsclr <= '0';
when s4022 => state := s4023; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4023 => 			--20
	if (addfprdy = '1') then state := s4024;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4023; end if;
when s4024 => state := s4025; 	--21
	addfpsclr <= '0';
when s4025 => state := s4026; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (238, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4026 => state := s4027; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (414, 12)); -- offset LSB 366
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s4027 => state := s4028;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (415, 12)); -- offset MSB 367
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4028 => state := s4029; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4029 => 			--4
	if (fixed2floatrdy = '1') then state := s4030;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4029; end if;
when s4030 => state := s4031; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4031 => 			--6
	if (mulfprdy = '1') then state := s4032;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4031; end if;
when s4032 => state := s4033; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4033 => 			--8
	if (mulfprdy = '1') then state := s4034;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4033; end if;
when s4034 => state := s4035; 	--9
	mulfpsclr <= '0';
when s4035 => state := s4036; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4036 => 			--11
	if (mulfprdy = '1') then state := s4037;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4036; end if;
when s4037 => state := s4038; 	--12
	mulfpsclr <= '0';
when s4038 => state := s4039; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4039 => 			--14
	if (addfprdy = '1') then state := s4040;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4039; end if;
when s4040 => state := s4041; 	--15
	addfpsclr <= '0';
when s4041 => state := s4042; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4042 => 			--17
	if (addfprdy = '1') then state := s4043;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4042; end if;
when s4043 => state := s4044; 	--18
	addfpsclr <= '0';
when s4044 => state := s4045; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4045 => 			--20
	if (addfprdy = '1') then state := s4046;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4045; end if;
when s4046 => state := s4047; 	--21
	addfpsclr <= '0';
when s4047 => state := s4048; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (239, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4048 => state := s4049; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (416, 12)); -- offset LSB 368
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s4049 => state := s4050;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (417, 12)); -- offset MSB 369
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4050 => state := s4051; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4051 => 			--4
	if (fixed2floatrdy = '1') then state := s4052;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4051; end if;
when s4052 => state := s4053; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4053 => 			--6
	if (mulfprdy = '1') then state := s4054;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4053; end if;
when s4054 => state := s4055; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4055 => 			--8
	if (mulfprdy = '1') then state := s4056;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4055; end if;
when s4056 => state := s4057; 	--9
	mulfpsclr <= '0';
when s4057 => state := s4058; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4058 => 			--11
	if (mulfprdy = '1') then state := s4059;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4058; end if;
when s4059 => state := s4060; 	--12
	mulfpsclr <= '0';
when s4060 => state := s4061; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4061 => 			--14
	if (addfprdy = '1') then state := s4062;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4061; end if;
when s4062 => state := s4063; 	--15
	addfpsclr <= '0';
when s4063 => state := s4064; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4064 => 			--17
	if (addfprdy = '1') then state := s4065;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4064; end if;
when s4065 => state := s4066; 	--18
	addfpsclr <= '0';
when s4066 => state := s4067; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4067 => 			--20
	if (addfprdy = '1') then state := s4068;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4067; end if;
when s4068 => state := s4069; 	--21
	addfpsclr <= '0';
when s4069 => state := s4070; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (240, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4070 => state := s4071; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (418, 12)); -- offset LSB 370
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s4071 => state := s4072;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (419, 12)); -- offset MSB 371
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4072 => state := s4073; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4073 => 			--4
	if (fixed2floatrdy = '1') then state := s4074;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4073; end if;
when s4074 => state := s4075; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4075 => 			--6
	if (mulfprdy = '1') then state := s4076;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4075; end if;
when s4076 => state := s4077; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4077 => 			--8
	if (mulfprdy = '1') then state := s4078;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4077; end if;
when s4078 => state := s4079; 	--9
	mulfpsclr <= '0';
when s4079 => state := s4080; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4080 => 			--11
	if (mulfprdy = '1') then state := s4081;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4080; end if;
when s4081 => state := s4082; 	--12
	mulfpsclr <= '0';
when s4082 => state := s4083; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4083 => 			--14
	if (addfprdy = '1') then state := s4084;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4083; end if;
when s4084 => state := s4085; 	--15
	addfpsclr <= '0';
when s4085 => state := s4086; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4086 => 			--17
	if (addfprdy = '1') then state := s4087;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4086; end if;
when s4087 => state := s4088; 	--18
	addfpsclr <= '0';
when s4088 => state := s4089; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4089 => 			--20
	if (addfprdy = '1') then state := s4090;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4089; end if;
when s4090 => state := s4091; 	--21
	addfpsclr <= '0';
when s4091 => state := s4092; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (241, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4092 => state := s4093; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (420, 12)); -- offset LSB 372
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s4093 => state := s4094;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (421, 12)); -- offset MSB 373
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4094 => state := s4095; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4095 => 			--4
	if (fixed2floatrdy = '1') then state := s4096;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4095; end if;
when s4096 => state := s4097; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4097 => 			--6
	if (mulfprdy = '1') then state := s4098;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4097; end if;
when s4098 => state := s4099; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4099 => 			--8
	if (mulfprdy = '1') then state := s4100;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4099; end if;
when s4100 => state := s4101; 	--9
	mulfpsclr <= '0';
when s4101 => state := s4102; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4102 => 			--11
	if (mulfprdy = '1') then state := s4103;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4102; end if;
when s4103 => state := s4104; 	--12
	mulfpsclr <= '0';
when s4104 => state := s4105; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4105 => 			--14
	if (addfprdy = '1') then state := s4106;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4105; end if;
when s4106 => state := s4107; 	--15
	addfpsclr <= '0';
when s4107 => state := s4108; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4108 => 			--17
	if (addfprdy = '1') then state := s4109;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4108; end if;
when s4109 => state := s4110; 	--18
	addfpsclr <= '0';
when s4110 => state := s4111; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4111 => 			--20
	if (addfprdy = '1') then state := s4112;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4111; end if;
when s4112 => state := s4113; 	--21
	addfpsclr <= '0';
when s4113 => state := s4114; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (242, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4114 => state := s4115; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (422, 12)); -- offset LSB 374
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s4115 => state := s4116;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (423, 12)); -- offset MSB 375
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4116 => state := s4117; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4117 => 			--4
	if (fixed2floatrdy = '1') then state := s4118;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4117; end if;
when s4118 => state := s4119; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4119 => 			--6
	if (mulfprdy = '1') then state := s4120;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4119; end if;
when s4120 => state := s4121; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4121 => 			--8
	if (mulfprdy = '1') then state := s4122;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4121; end if;
when s4122 => state := s4123; 	--9
	mulfpsclr <= '0';
when s4123 => state := s4124; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4124 => 			--11
	if (mulfprdy = '1') then state := s4125;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4124; end if;
when s4125 => state := s4126; 	--12
	mulfpsclr <= '0';
when s4126 => state := s4127; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4127 => 			--14
	if (addfprdy = '1') then state := s4128;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4127; end if;
when s4128 => state := s4129; 	--15
	addfpsclr <= '0';
when s4129 => state := s4130; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4130 => 			--17
	if (addfprdy = '1') then state := s4131;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4130; end if;
when s4131 => state := s4132; 	--18
	addfpsclr <= '0';
when s4132 => state := s4133; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4133 => 			--20
	if (addfprdy = '1') then state := s4134;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4133; end if;
when s4134 => state := s4135; 	--21
	addfpsclr <= '0';
when s4135 => state := s4136; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (243, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4136 => state := s4137; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (424, 12)); -- offset LSB 376
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s4137 => state := s4138;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (425, 12)); -- offset MSB 377
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4138 => state := s4139; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4139 => 			--4
	if (fixed2floatrdy = '1') then state := s4140;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4139; end if;
when s4140 => state := s4141; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4141 => 			--6
	if (mulfprdy = '1') then state := s4142;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4141; end if;
when s4142 => state := s4143; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4143 => 			--8
	if (mulfprdy = '1') then state := s4144;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4143; end if;
when s4144 => state := s4145; 	--9
	mulfpsclr <= '0';
when s4145 => state := s4146; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4146 => 			--11
	if (mulfprdy = '1') then state := s4147;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4146; end if;
when s4147 => state := s4148; 	--12
	mulfpsclr <= '0';
when s4148 => state := s4149; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4149 => 			--14
	if (addfprdy = '1') then state := s4150;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4149; end if;
when s4150 => state := s4151; 	--15
	addfpsclr <= '0';
when s4151 => state := s4152; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4152 => 			--17
	if (addfprdy = '1') then state := s4153;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4152; end if;
when s4153 => state := s4154; 	--18
	addfpsclr <= '0';
when s4154 => state := s4155; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4155 => 			--20
	if (addfprdy = '1') then state := s4156;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4155; end if;
when s4156 => state := s4157; 	--21
	addfpsclr <= '0';
when s4157 => state := s4158; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (244, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4158 => state := s4159; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (426, 12)); -- offset LSB 378
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s4159 => state := s4160;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (427, 12)); -- offset MSB 379
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4160 => state := s4161; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4161 => 			--4
	if (fixed2floatrdy = '1') then state := s4162;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4161; end if;
when s4162 => state := s4163; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4163 => 			--6
	if (mulfprdy = '1') then state := s4164;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4163; end if;
when s4164 => state := s4165; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4165 => 			--8
	if (mulfprdy = '1') then state := s4166;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4165; end if;
when s4166 => state := s4167; 	--9
	mulfpsclr <= '0';
when s4167 => state := s4168; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4168 => 			--11
	if (mulfprdy = '1') then state := s4169;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4168; end if;
when s4169 => state := s4170; 	--12
	mulfpsclr <= '0';
when s4170 => state := s4171; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4171 => 			--14
	if (addfprdy = '1') then state := s4172;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4171; end if;
when s4172 => state := s4173; 	--15
	addfpsclr <= '0';
when s4173 => state := s4174; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4174 => 			--17
	if (addfprdy = '1') then state := s4175;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4174; end if;
when s4175 => state := s4176; 	--18
	addfpsclr <= '0';
when s4176 => state := s4177; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4177 => 			--20
	if (addfprdy = '1') then state := s4178;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4177; end if;
when s4178 => state := s4179; 	--21
	addfpsclr <= '0';
when s4179 => state := s4180; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (245, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4180 => state := s4181; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (428, 12)); -- offset LSB 380
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s4181 => state := s4182;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (429, 12)); -- offset MSB 381
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4182 => state := s4183; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4183 => 			--4
	if (fixed2floatrdy = '1') then state := s4184;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4183; end if;
when s4184 => state := s4185; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4185 => 			--6
	if (mulfprdy = '1') then state := s4186;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4185; end if;
when s4186 => state := s4187; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4187 => 			--8
	if (mulfprdy = '1') then state := s4188;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4187; end if;
when s4188 => state := s4189; 	--9
	mulfpsclr <= '0';
when s4189 => state := s4190; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4190 => 			--11
	if (mulfprdy = '1') then state := s4191;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4190; end if;
when s4191 => state := s4192; 	--12
	mulfpsclr <= '0';
when s4192 => state := s4193; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4193 => 			--14
	if (addfprdy = '1') then state := s4194;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4193; end if;
when s4194 => state := s4195; 	--15
	addfpsclr <= '0';
when s4195 => state := s4196; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4196 => 			--17
	if (addfprdy = '1') then state := s4197;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4196; end if;
when s4197 => state := s4198; 	--18
	addfpsclr <= '0';
when s4198 => state := s4199; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4199 => 			--20
	if (addfprdy = '1') then state := s4200;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4199; end if;
when s4200 => state := s4201; 	--21
	addfpsclr <= '0';
when s4201 => state := s4202; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (246, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4202 => state := s4203; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (430, 12)); -- offset LSB 382
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s4203 => state := s4204;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (431, 12)); -- offset MSB 383
	addra <= std_logic_vector (to_unsigned (5, 10)); -- OCCrowI 5
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4204 => state := s4205; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4205 => 			--4
	if (fixed2floatrdy = '1') then state := s4206;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4205; end if;
when s4206 => state := s4207; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4207 => 			--6
	if (mulfprdy = '1') then state := s4208;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4207; end if;
when s4208 => state := s4209; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4209 => 			--8
	if (mulfprdy = '1') then state := s4210;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4209; end if;
when s4210 => state := s4211; 	--9
	mulfpsclr <= '0';
when s4211 => state := s4212; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4212 => 			--11
	if (mulfprdy = '1') then state := s4213;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4212; end if;
when s4213 => state := s4214; 	--12
	mulfpsclr <= '0';
when s4214 => state := s4215; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4215 => 			--14
	if (addfprdy = '1') then state := s4216;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4215; end if;
when s4216 => state := s4217; 	--15
	addfpsclr <= '0';
when s4217 => state := s4218; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4218 => 			--17
	if (addfprdy = '1') then state := s4219;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4218; end if;
when s4219 => state := s4220; 	--18
	addfpsclr <= '0';
when s4220 => state := s4221; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4221 => 			--20
	if (addfprdy = '1') then state := s4222;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4221; end if;
when s4222 => state := s4223; 	--21
	addfpsclr <= '0';
when s4223 => state := s4224; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (247, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4224 => state := s4225; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (432, 12)); -- offset LSB 384
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s4225 => state := s4226;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (433, 12)); -- offset MSB 385
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4226 => state := s4227; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4227 => 			--4
	if (fixed2floatrdy = '1') then state := s4228;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4227; end if;
when s4228 => state := s4229; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4229 => 			--6
	if (mulfprdy = '1') then state := s4230;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4229; end if;
when s4230 => state := s4231; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4231 => 			--8
	if (mulfprdy = '1') then state := s4232;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4231; end if;
when s4232 => state := s4233; 	--9
	mulfpsclr <= '0';
when s4233 => state := s4234; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4234 => 			--11
	if (mulfprdy = '1') then state := s4235;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4234; end if;
when s4235 => state := s4236; 	--12
	mulfpsclr <= '0';
when s4236 => state := s4237; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4237 => 			--14
	if (addfprdy = '1') then state := s4238;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4237; end if;
when s4238 => state := s4239; 	--15
	addfpsclr <= '0';
when s4239 => state := s4240; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4240 => 			--17
	if (addfprdy = '1') then state := s4241;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4240; end if;
when s4241 => state := s4242; 	--18
	addfpsclr <= '0';
when s4242 => state := s4243; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4243 => 			--20
	if (addfprdy = '1') then state := s4244;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4243; end if;
when s4244 => state := s4245; 	--21
	addfpsclr <= '0';
when s4245 => state := s4246; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (248, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4246 => state := s4247; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (434, 12)); -- offset LSB 386
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s4247 => state := s4248;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (435, 12)); -- offset MSB 387
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4248 => state := s4249; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4249 => 			--4
	if (fixed2floatrdy = '1') then state := s4250;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4249; end if;
when s4250 => state := s4251; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4251 => 			--6
	if (mulfprdy = '1') then state := s4252;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4251; end if;
when s4252 => state := s4253; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4253 => 			--8
	if (mulfprdy = '1') then state := s4254;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4253; end if;
when s4254 => state := s4255; 	--9
	mulfpsclr <= '0';
when s4255 => state := s4256; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4256 => 			--11
	if (mulfprdy = '1') then state := s4257;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4256; end if;
when s4257 => state := s4258; 	--12
	mulfpsclr <= '0';
when s4258 => state := s4259; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4259 => 			--14
	if (addfprdy = '1') then state := s4260;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4259; end if;
when s4260 => state := s4261; 	--15
	addfpsclr <= '0';
when s4261 => state := s4262; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4262 => 			--17
	if (addfprdy = '1') then state := s4263;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4262; end if;
when s4263 => state := s4264; 	--18
	addfpsclr <= '0';
when s4264 => state := s4265; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4265 => 			--20
	if (addfprdy = '1') then state := s4266;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4265; end if;
when s4266 => state := s4267; 	--21
	addfpsclr <= '0';
when s4267 => state := s4268; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (249, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4268 => state := s4269; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (436, 12)); -- offset LSB 388
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s4269 => state := s4270;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (437, 12)); -- offset MSB 389
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4270 => state := s4271; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4271 => 			--4
	if (fixed2floatrdy = '1') then state := s4272;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4271; end if;
when s4272 => state := s4273; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4273 => 			--6
	if (mulfprdy = '1') then state := s4274;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4273; end if;
when s4274 => state := s4275; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4275 => 			--8
	if (mulfprdy = '1') then state := s4276;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4275; end if;
when s4276 => state := s4277; 	--9
	mulfpsclr <= '0';
when s4277 => state := s4278; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4278 => 			--11
	if (mulfprdy = '1') then state := s4279;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4278; end if;
when s4279 => state := s4280; 	--12
	mulfpsclr <= '0';
when s4280 => state := s4281; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4281 => 			--14
	if (addfprdy = '1') then state := s4282;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4281; end if;
when s4282 => state := s4283; 	--15
	addfpsclr <= '0';
when s4283 => state := s4284; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4284 => 			--17
	if (addfprdy = '1') then state := s4285;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4284; end if;
when s4285 => state := s4286; 	--18
	addfpsclr <= '0';
when s4286 => state := s4287; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4287 => 			--20
	if (addfprdy = '1') then state := s4288;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4287; end if;
when s4288 => state := s4289; 	--21
	addfpsclr <= '0';
when s4289 => state := s4290; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (250, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4290 => state := s4291; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (438, 12)); -- offset LSB 390
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s4291 => state := s4292;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (439, 12)); -- offset MSB 391
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4292 => state := s4293; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4293 => 			--4
	if (fixed2floatrdy = '1') then state := s4294;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4293; end if;
when s4294 => state := s4295; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4295 => 			--6
	if (mulfprdy = '1') then state := s4296;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4295; end if;
when s4296 => state := s4297; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4297 => 			--8
	if (mulfprdy = '1') then state := s4298;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4297; end if;
when s4298 => state := s4299; 	--9
	mulfpsclr <= '0';
when s4299 => state := s4300; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4300 => 			--11
	if (mulfprdy = '1') then state := s4301;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4300; end if;
when s4301 => state := s4302; 	--12
	mulfpsclr <= '0';
when s4302 => state := s4303; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4303 => 			--14
	if (addfprdy = '1') then state := s4304;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4303; end if;
when s4304 => state := s4305; 	--15
	addfpsclr <= '0';
when s4305 => state := s4306; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4306 => 			--17
	if (addfprdy = '1') then state := s4307;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4306; end if;
when s4307 => state := s4308; 	--18
	addfpsclr <= '0';
when s4308 => state := s4309; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4309 => 			--20
	if (addfprdy = '1') then state := s4310;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4309; end if;
when s4310 => state := s4311; 	--21
	addfpsclr <= '0';
when s4311 => state := s4312; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (251, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4312 => state := s4313; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (440, 12)); -- offset LSB 392
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s4313 => state := s4314;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (441, 12)); -- offset MSB 393
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4314 => state := s4315; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4315 => 			--4
	if (fixed2floatrdy = '1') then state := s4316;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4315; end if;
when s4316 => state := s4317; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4317 => 			--6
	if (mulfprdy = '1') then state := s4318;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4317; end if;
when s4318 => state := s4319; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4319 => 			--8
	if (mulfprdy = '1') then state := s4320;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4319; end if;
when s4320 => state := s4321; 	--9
	mulfpsclr <= '0';
when s4321 => state := s4322; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4322 => 			--11
	if (mulfprdy = '1') then state := s4323;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4322; end if;
when s4323 => state := s4324; 	--12
	mulfpsclr <= '0';
when s4324 => state := s4325; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4325 => 			--14
	if (addfprdy = '1') then state := s4326;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4325; end if;
when s4326 => state := s4327; 	--15
	addfpsclr <= '0';
when s4327 => state := s4328; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4328 => 			--17
	if (addfprdy = '1') then state := s4329;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4328; end if;
when s4329 => state := s4330; 	--18
	addfpsclr <= '0';
when s4330 => state := s4331; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4331 => 			--20
	if (addfprdy = '1') then state := s4332;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4331; end if;
when s4332 => state := s4333; 	--21
	addfpsclr <= '0';
when s4333 => state := s4334; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (252, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4334 => state := s4335; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (442, 12)); -- offset LSB 394
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s4335 => state := s4336;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (443, 12)); -- offset MSB 395
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4336 => state := s4337; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4337 => 			--4
	if (fixed2floatrdy = '1') then state := s4338;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4337; end if;
when s4338 => state := s4339; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4339 => 			--6
	if (mulfprdy = '1') then state := s4340;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4339; end if;
when s4340 => state := s4341; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4341 => 			--8
	if (mulfprdy = '1') then state := s4342;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4341; end if;
when s4342 => state := s4343; 	--9
	mulfpsclr <= '0';
when s4343 => state := s4344; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4344 => 			--11
	if (mulfprdy = '1') then state := s4345;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4344; end if;
when s4345 => state := s4346; 	--12
	mulfpsclr <= '0';
when s4346 => state := s4347; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4347 => 			--14
	if (addfprdy = '1') then state := s4348;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4347; end if;
when s4348 => state := s4349; 	--15
	addfpsclr <= '0';
when s4349 => state := s4350; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4350 => 			--17
	if (addfprdy = '1') then state := s4351;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4350; end if;
when s4351 => state := s4352; 	--18
	addfpsclr <= '0';
when s4352 => state := s4353; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4353 => 			--20
	if (addfprdy = '1') then state := s4354;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4353; end if;
when s4354 => state := s4355; 	--21
	addfpsclr <= '0';
when s4355 => state := s4356; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (253, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4356 => state := s4357; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (444, 12)); -- offset LSB 396
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s4357 => state := s4358;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (445, 12)); -- offset MSB 397
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4358 => state := s4359; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4359 => 			--4
	if (fixed2floatrdy = '1') then state := s4360;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4359; end if;
when s4360 => state := s4361; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4361 => 			--6
	if (mulfprdy = '1') then state := s4362;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4361; end if;
when s4362 => state := s4363; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4363 => 			--8
	if (mulfprdy = '1') then state := s4364;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4363; end if;
when s4364 => state := s4365; 	--9
	mulfpsclr <= '0';
when s4365 => state := s4366; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4366 => 			--11
	if (mulfprdy = '1') then state := s4367;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4366; end if;
when s4367 => state := s4368; 	--12
	mulfpsclr <= '0';
when s4368 => state := s4369; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4369 => 			--14
	if (addfprdy = '1') then state := s4370;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4369; end if;
when s4370 => state := s4371; 	--15
	addfpsclr <= '0';
when s4371 => state := s4372; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4372 => 			--17
	if (addfprdy = '1') then state := s4373;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4372; end if;
when s4373 => state := s4374; 	--18
	addfpsclr <= '0';
when s4374 => state := s4375; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4375 => 			--20
	if (addfprdy = '1') then state := s4376;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4375; end if;
when s4376 => state := s4377; 	--21
	addfpsclr <= '0';
when s4377 => state := s4378; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (254, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4378 => state := s4379; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (446, 12)); -- offset LSB 398
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s4379 => state := s4380;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (447, 12)); -- offset MSB 399
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4380 => state := s4381; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4381 => 			--4
	if (fixed2floatrdy = '1') then state := s4382;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4381; end if;
when s4382 => state := s4383; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4383 => 			--6
	if (mulfprdy = '1') then state := s4384;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4383; end if;
when s4384 => state := s4385; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4385 => 			--8
	if (mulfprdy = '1') then state := s4386;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4385; end if;
when s4386 => state := s4387; 	--9
	mulfpsclr <= '0';
when s4387 => state := s4388; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4388 => 			--11
	if (mulfprdy = '1') then state := s4389;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4388; end if;
when s4389 => state := s4390; 	--12
	mulfpsclr <= '0';
when s4390 => state := s4391; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4391 => 			--14
	if (addfprdy = '1') then state := s4392;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4391; end if;
when s4392 => state := s4393; 	--15
	addfpsclr <= '0';
when s4393 => state := s4394; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4394 => 			--17
	if (addfprdy = '1') then state := s4395;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4394; end if;
when s4395 => state := s4396; 	--18
	addfpsclr <= '0';
when s4396 => state := s4397; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4397 => 			--20
	if (addfprdy = '1') then state := s4398;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4397; end if;
when s4398 => state := s4399; 	--21
	addfpsclr <= '0';
when s4399 => state := s4400; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (255, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4400 => state := s4401; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (448, 12)); -- offset LSB 400
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s4401 => state := s4402;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (449, 12)); -- offset MSB 401
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4402 => state := s4403; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4403 => 			--4
	if (fixed2floatrdy = '1') then state := s4404;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4403; end if;
when s4404 => state := s4405; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4405 => 			--6
	if (mulfprdy = '1') then state := s4406;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4405; end if;
when s4406 => state := s4407; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4407 => 			--8
	if (mulfprdy = '1') then state := s4408;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4407; end if;
when s4408 => state := s4409; 	--9
	mulfpsclr <= '0';
when s4409 => state := s4410; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4410 => 			--11
	if (mulfprdy = '1') then state := s4411;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4410; end if;
when s4411 => state := s4412; 	--12
	mulfpsclr <= '0';
when s4412 => state := s4413; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4413 => 			--14
	if (addfprdy = '1') then state := s4414;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4413; end if;
when s4414 => state := s4415; 	--15
	addfpsclr <= '0';
when s4415 => state := s4416; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4416 => 			--17
	if (addfprdy = '1') then state := s4417;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4416; end if;
when s4417 => state := s4418; 	--18
	addfpsclr <= '0';
when s4418 => state := s4419; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4419 => 			--20
	if (addfprdy = '1') then state := s4420;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4419; end if;
when s4420 => state := s4421; 	--21
	addfpsclr <= '0';
when s4421 => state := s4422; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (256, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4422 => state := s4423; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (450, 12)); -- offset LSB 402
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s4423 => state := s4424;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (451, 12)); -- offset MSB 403
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4424 => state := s4425; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4425 => 			--4
	if (fixed2floatrdy = '1') then state := s4426;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4425; end if;
when s4426 => state := s4427; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4427 => 			--6
	if (mulfprdy = '1') then state := s4428;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4427; end if;
when s4428 => state := s4429; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4429 => 			--8
	if (mulfprdy = '1') then state := s4430;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4429; end if;
when s4430 => state := s4431; 	--9
	mulfpsclr <= '0';
when s4431 => state := s4432; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4432 => 			--11
	if (mulfprdy = '1') then state := s4433;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4432; end if;
when s4433 => state := s4434; 	--12
	mulfpsclr <= '0';
when s4434 => state := s4435; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4435 => 			--14
	if (addfprdy = '1') then state := s4436;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4435; end if;
when s4436 => state := s4437; 	--15
	addfpsclr <= '0';
when s4437 => state := s4438; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4438 => 			--17
	if (addfprdy = '1') then state := s4439;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4438; end if;
when s4439 => state := s4440; 	--18
	addfpsclr <= '0';
when s4440 => state := s4441; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4441 => 			--20
	if (addfprdy = '1') then state := s4442;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4441; end if;
when s4442 => state := s4443; 	--21
	addfpsclr <= '0';
when s4443 => state := s4444; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (257, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4444 => state := s4445; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (452, 12)); -- offset LSB 404
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s4445 => state := s4446;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (453, 12)); -- offset MSB 405
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4446 => state := s4447; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4447 => 			--4
	if (fixed2floatrdy = '1') then state := s4448;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4447; end if;
when s4448 => state := s4449; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4449 => 			--6
	if (mulfprdy = '1') then state := s4450;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4449; end if;
when s4450 => state := s4451; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4451 => 			--8
	if (mulfprdy = '1') then state := s4452;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4451; end if;
when s4452 => state := s4453; 	--9
	mulfpsclr <= '0';
when s4453 => state := s4454; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4454 => 			--11
	if (mulfprdy = '1') then state := s4455;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4454; end if;
when s4455 => state := s4456; 	--12
	mulfpsclr <= '0';
when s4456 => state := s4457; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4457 => 			--14
	if (addfprdy = '1') then state := s4458;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4457; end if;
when s4458 => state := s4459; 	--15
	addfpsclr <= '0';
when s4459 => state := s4460; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4460 => 			--17
	if (addfprdy = '1') then state := s4461;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4460; end if;
when s4461 => state := s4462; 	--18
	addfpsclr <= '0';
when s4462 => state := s4463; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4463 => 			--20
	if (addfprdy = '1') then state := s4464;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4463; end if;
when s4464 => state := s4465; 	--21
	addfpsclr <= '0';
when s4465 => state := s4466; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (258, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4466 => state := s4467; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (454, 12)); -- offset LSB 406
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s4467 => state := s4468;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (455, 12)); -- offset MSB 407
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4468 => state := s4469; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4469 => 			--4
	if (fixed2floatrdy = '1') then state := s4470;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4469; end if;
when s4470 => state := s4471; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4471 => 			--6
	if (mulfprdy = '1') then state := s4472;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4471; end if;
when s4472 => state := s4473; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4473 => 			--8
	if (mulfprdy = '1') then state := s4474;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4473; end if;
when s4474 => state := s4475; 	--9
	mulfpsclr <= '0';
when s4475 => state := s4476; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4476 => 			--11
	if (mulfprdy = '1') then state := s4477;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4476; end if;
when s4477 => state := s4478; 	--12
	mulfpsclr <= '0';
when s4478 => state := s4479; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4479 => 			--14
	if (addfprdy = '1') then state := s4480;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4479; end if;
when s4480 => state := s4481; 	--15
	addfpsclr <= '0';
when s4481 => state := s4482; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4482 => 			--17
	if (addfprdy = '1') then state := s4483;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4482; end if;
when s4483 => state := s4484; 	--18
	addfpsclr <= '0';
when s4484 => state := s4485; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4485 => 			--20
	if (addfprdy = '1') then state := s4486;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4485; end if;
when s4486 => state := s4487; 	--21
	addfpsclr <= '0';
when s4487 => state := s4488; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (259, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4488 => state := s4489; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (456, 12)); -- offset LSB 408
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s4489 => state := s4490;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (457, 12)); -- offset MSB 409
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4490 => state := s4491; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4491 => 			--4
	if (fixed2floatrdy = '1') then state := s4492;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4491; end if;
when s4492 => state := s4493; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4493 => 			--6
	if (mulfprdy = '1') then state := s4494;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4493; end if;
when s4494 => state := s4495; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4495 => 			--8
	if (mulfprdy = '1') then state := s4496;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4495; end if;
when s4496 => state := s4497; 	--9
	mulfpsclr <= '0';
when s4497 => state := s4498; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4498 => 			--11
	if (mulfprdy = '1') then state := s4499;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4498; end if;
when s4499 => state := s4500; 	--12
	mulfpsclr <= '0';
when s4500 => state := s4501; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4501 => 			--14
	if (addfprdy = '1') then state := s4502;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4501; end if;
when s4502 => state := s4503; 	--15
	addfpsclr <= '0';
when s4503 => state := s4504; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4504 => 			--17
	if (addfprdy = '1') then state := s4505;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4504; end if;
when s4505 => state := s4506; 	--18
	addfpsclr <= '0';
when s4506 => state := s4507; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4507 => 			--20
	if (addfprdy = '1') then state := s4508;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4507; end if;
when s4508 => state := s4509; 	--21
	addfpsclr <= '0';
when s4509 => state := s4510; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (260, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4510 => state := s4511; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (458, 12)); -- offset LSB 410
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s4511 => state := s4512;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (459, 12)); -- offset MSB 411
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4512 => state := s4513; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4513 => 			--4
	if (fixed2floatrdy = '1') then state := s4514;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4513; end if;
when s4514 => state := s4515; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4515 => 			--6
	if (mulfprdy = '1') then state := s4516;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4515; end if;
when s4516 => state := s4517; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4517 => 			--8
	if (mulfprdy = '1') then state := s4518;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4517; end if;
when s4518 => state := s4519; 	--9
	mulfpsclr <= '0';
when s4519 => state := s4520; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4520 => 			--11
	if (mulfprdy = '1') then state := s4521;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4520; end if;
when s4521 => state := s4522; 	--12
	mulfpsclr <= '0';
when s4522 => state := s4523; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4523 => 			--14
	if (addfprdy = '1') then state := s4524;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4523; end if;
when s4524 => state := s4525; 	--15
	addfpsclr <= '0';
when s4525 => state := s4526; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4526 => 			--17
	if (addfprdy = '1') then state := s4527;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4526; end if;
when s4527 => state := s4528; 	--18
	addfpsclr <= '0';
when s4528 => state := s4529; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4529 => 			--20
	if (addfprdy = '1') then state := s4530;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4529; end if;
when s4530 => state := s4531; 	--21
	addfpsclr <= '0';
when s4531 => state := s4532; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (261, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4532 => state := s4533; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (460, 12)); -- offset LSB 412
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s4533 => state := s4534;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (461, 12)); -- offset MSB 413
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4534 => state := s4535; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4535 => 			--4
	if (fixed2floatrdy = '1') then state := s4536;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4535; end if;
when s4536 => state := s4537; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4537 => 			--6
	if (mulfprdy = '1') then state := s4538;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4537; end if;
when s4538 => state := s4539; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4539 => 			--8
	if (mulfprdy = '1') then state := s4540;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4539; end if;
when s4540 => state := s4541; 	--9
	mulfpsclr <= '0';
when s4541 => state := s4542; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4542 => 			--11
	if (mulfprdy = '1') then state := s4543;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4542; end if;
when s4543 => state := s4544; 	--12
	mulfpsclr <= '0';
when s4544 => state := s4545; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4545 => 			--14
	if (addfprdy = '1') then state := s4546;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4545; end if;
when s4546 => state := s4547; 	--15
	addfpsclr <= '0';
when s4547 => state := s4548; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4548 => 			--17
	if (addfprdy = '1') then state := s4549;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4548; end if;
when s4549 => state := s4550; 	--18
	addfpsclr <= '0';
when s4550 => state := s4551; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4551 => 			--20
	if (addfprdy = '1') then state := s4552;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4551; end if;
when s4552 => state := s4553; 	--21
	addfpsclr <= '0';
when s4553 => state := s4554; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (262, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4554 => state := s4555; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (462, 12)); -- offset LSB 414
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s4555 => state := s4556;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (463, 12)); -- offset MSB 415
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4556 => state := s4557; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4557 => 			--4
	if (fixed2floatrdy = '1') then state := s4558;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4557; end if;
when s4558 => state := s4559; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4559 => 			--6
	if (mulfprdy = '1') then state := s4560;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4559; end if;
when s4560 => state := s4561; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4561 => 			--8
	if (mulfprdy = '1') then state := s4562;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4561; end if;
when s4562 => state := s4563; 	--9
	mulfpsclr <= '0';
when s4563 => state := s4564; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4564 => 			--11
	if (mulfprdy = '1') then state := s4565;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4564; end if;
when s4565 => state := s4566; 	--12
	mulfpsclr <= '0';
when s4566 => state := s4567; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4567 => 			--14
	if (addfprdy = '1') then state := s4568;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4567; end if;
when s4568 => state := s4569; 	--15
	addfpsclr <= '0';
when s4569 => state := s4570; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4570 => 			--17
	if (addfprdy = '1') then state := s4571;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4570; end if;
when s4571 => state := s4572; 	--18
	addfpsclr <= '0';
when s4572 => state := s4573; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4573 => 			--20
	if (addfprdy = '1') then state := s4574;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4573; end if;
when s4574 => state := s4575; 	--21
	addfpsclr <= '0';
when s4575 => state := s4576; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (263, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4576 => state := s4577; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (464, 12)); -- offset LSB 416
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s4577 => state := s4578;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (465, 12)); -- offset MSB 417
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4578 => state := s4579; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4579 => 			--4
	if (fixed2floatrdy = '1') then state := s4580;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4579; end if;
when s4580 => state := s4581; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4581 => 			--6
	if (mulfprdy = '1') then state := s4582;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4581; end if;
when s4582 => state := s4583; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4583 => 			--8
	if (mulfprdy = '1') then state := s4584;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4583; end if;
when s4584 => state := s4585; 	--9
	mulfpsclr <= '0';
when s4585 => state := s4586; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4586 => 			--11
	if (mulfprdy = '1') then state := s4587;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4586; end if;
when s4587 => state := s4588; 	--12
	mulfpsclr <= '0';
when s4588 => state := s4589; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4589 => 			--14
	if (addfprdy = '1') then state := s4590;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4589; end if;
when s4590 => state := s4591; 	--15
	addfpsclr <= '0';
when s4591 => state := s4592; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4592 => 			--17
	if (addfprdy = '1') then state := s4593;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4592; end if;
when s4593 => state := s4594; 	--18
	addfpsclr <= '0';
when s4594 => state := s4595; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4595 => 			--20
	if (addfprdy = '1') then state := s4596;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4595; end if;
when s4596 => state := s4597; 	--21
	addfpsclr <= '0';
when s4597 => state := s4598; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (264, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4598 => state := s4599; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (466, 12)); -- offset LSB 418
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s4599 => state := s4600;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (467, 12)); -- offset MSB 419
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4600 => state := s4601; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4601 => 			--4
	if (fixed2floatrdy = '1') then state := s4602;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4601; end if;
when s4602 => state := s4603; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4603 => 			--6
	if (mulfprdy = '1') then state := s4604;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4603; end if;
when s4604 => state := s4605; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4605 => 			--8
	if (mulfprdy = '1') then state := s4606;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4605; end if;
when s4606 => state := s4607; 	--9
	mulfpsclr <= '0';
when s4607 => state := s4608; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4608 => 			--11
	if (mulfprdy = '1') then state := s4609;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4608; end if;
when s4609 => state := s4610; 	--12
	mulfpsclr <= '0';
when s4610 => state := s4611; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4611 => 			--14
	if (addfprdy = '1') then state := s4612;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4611; end if;
when s4612 => state := s4613; 	--15
	addfpsclr <= '0';
when s4613 => state := s4614; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4614 => 			--17
	if (addfprdy = '1') then state := s4615;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4614; end if;
when s4615 => state := s4616; 	--18
	addfpsclr <= '0';
when s4616 => state := s4617; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4617 => 			--20
	if (addfprdy = '1') then state := s4618;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4617; end if;
when s4618 => state := s4619; 	--21
	addfpsclr <= '0';
when s4619 => state := s4620; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (265, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4620 => state := s4621; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (468, 12)); -- offset LSB 420
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s4621 => state := s4622;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (469, 12)); -- offset MSB 421
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4622 => state := s4623; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4623 => 			--4
	if (fixed2floatrdy = '1') then state := s4624;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4623; end if;
when s4624 => state := s4625; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4625 => 			--6
	if (mulfprdy = '1') then state := s4626;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4625; end if;
when s4626 => state := s4627; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4627 => 			--8
	if (mulfprdy = '1') then state := s4628;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4627; end if;
when s4628 => state := s4629; 	--9
	mulfpsclr <= '0';
when s4629 => state := s4630; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4630 => 			--11
	if (mulfprdy = '1') then state := s4631;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4630; end if;
when s4631 => state := s4632; 	--12
	mulfpsclr <= '0';
when s4632 => state := s4633; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4633 => 			--14
	if (addfprdy = '1') then state := s4634;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4633; end if;
when s4634 => state := s4635; 	--15
	addfpsclr <= '0';
when s4635 => state := s4636; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4636 => 			--17
	if (addfprdy = '1') then state := s4637;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4636; end if;
when s4637 => state := s4638; 	--18
	addfpsclr <= '0';
when s4638 => state := s4639; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4639 => 			--20
	if (addfprdy = '1') then state := s4640;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4639; end if;
when s4640 => state := s4641; 	--21
	addfpsclr <= '0';
when s4641 => state := s4642; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (266, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4642 => state := s4643; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (470, 12)); -- offset LSB 422
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s4643 => state := s4644;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (471, 12)); -- offset MSB 423
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4644 => state := s4645; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4645 => 			--4
	if (fixed2floatrdy = '1') then state := s4646;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4645; end if;
when s4646 => state := s4647; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4647 => 			--6
	if (mulfprdy = '1') then state := s4648;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4647; end if;
when s4648 => state := s4649; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4649 => 			--8
	if (mulfprdy = '1') then state := s4650;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4649; end if;
when s4650 => state := s4651; 	--9
	mulfpsclr <= '0';
when s4651 => state := s4652; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4652 => 			--11
	if (mulfprdy = '1') then state := s4653;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4652; end if;
when s4653 => state := s4654; 	--12
	mulfpsclr <= '0';
when s4654 => state := s4655; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4655 => 			--14
	if (addfprdy = '1') then state := s4656;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4655; end if;
when s4656 => state := s4657; 	--15
	addfpsclr <= '0';
when s4657 => state := s4658; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4658 => 			--17
	if (addfprdy = '1') then state := s4659;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4658; end if;
when s4659 => state := s4660; 	--18
	addfpsclr <= '0';
when s4660 => state := s4661; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4661 => 			--20
	if (addfprdy = '1') then state := s4662;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4661; end if;
when s4662 => state := s4663; 	--21
	addfpsclr <= '0';
when s4663 => state := s4664; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (267, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4664 => state := s4665; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (472, 12)); -- offset LSB 424
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s4665 => state := s4666;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (473, 12)); -- offset MSB 425
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4666 => state := s4667; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4667 => 			--4
	if (fixed2floatrdy = '1') then state := s4668;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4667; end if;
when s4668 => state := s4669; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4669 => 			--6
	if (mulfprdy = '1') then state := s4670;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4669; end if;
when s4670 => state := s4671; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4671 => 			--8
	if (mulfprdy = '1') then state := s4672;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4671; end if;
when s4672 => state := s4673; 	--9
	mulfpsclr <= '0';
when s4673 => state := s4674; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4674 => 			--11
	if (mulfprdy = '1') then state := s4675;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4674; end if;
when s4675 => state := s4676; 	--12
	mulfpsclr <= '0';
when s4676 => state := s4677; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4677 => 			--14
	if (addfprdy = '1') then state := s4678;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4677; end if;
when s4678 => state := s4679; 	--15
	addfpsclr <= '0';
when s4679 => state := s4680; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4680 => 			--17
	if (addfprdy = '1') then state := s4681;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4680; end if;
when s4681 => state := s4682; 	--18
	addfpsclr <= '0';
when s4682 => state := s4683; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4683 => 			--20
	if (addfprdy = '1') then state := s4684;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4683; end if;
when s4684 => state := s4685; 	--21
	addfpsclr <= '0';
when s4685 => state := s4686; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (268, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4686 => state := s4687; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (474, 12)); -- offset LSB 426
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s4687 => state := s4688;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (475, 12)); -- offset MSB 427
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4688 => state := s4689; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4689 => 			--4
	if (fixed2floatrdy = '1') then state := s4690;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4689; end if;
when s4690 => state := s4691; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4691 => 			--6
	if (mulfprdy = '1') then state := s4692;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4691; end if;
when s4692 => state := s4693; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4693 => 			--8
	if (mulfprdy = '1') then state := s4694;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4693; end if;
when s4694 => state := s4695; 	--9
	mulfpsclr <= '0';
when s4695 => state := s4696; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4696 => 			--11
	if (mulfprdy = '1') then state := s4697;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4696; end if;
when s4697 => state := s4698; 	--12
	mulfpsclr <= '0';
when s4698 => state := s4699; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4699 => 			--14
	if (addfprdy = '1') then state := s4700;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4699; end if;
when s4700 => state := s4701; 	--15
	addfpsclr <= '0';
when s4701 => state := s4702; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4702 => 			--17
	if (addfprdy = '1') then state := s4703;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4702; end if;
when s4703 => state := s4704; 	--18
	addfpsclr <= '0';
when s4704 => state := s4705; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4705 => 			--20
	if (addfprdy = '1') then state := s4706;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4705; end if;
when s4706 => state := s4707; 	--21
	addfpsclr <= '0';
when s4707 => state := s4708; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (269, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4708 => state := s4709; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (476, 12)); -- offset LSB 428
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s4709 => state := s4710;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (477, 12)); -- offset MSB 429
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4710 => state := s4711; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4711 => 			--4
	if (fixed2floatrdy = '1') then state := s4712;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4711; end if;
when s4712 => state := s4713; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4713 => 			--6
	if (mulfprdy = '1') then state := s4714;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4713; end if;
when s4714 => state := s4715; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4715 => 			--8
	if (mulfprdy = '1') then state := s4716;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4715; end if;
when s4716 => state := s4717; 	--9
	mulfpsclr <= '0';
when s4717 => state := s4718; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4718 => 			--11
	if (mulfprdy = '1') then state := s4719;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4718; end if;
when s4719 => state := s4720; 	--12
	mulfpsclr <= '0';
when s4720 => state := s4721; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4721 => 			--14
	if (addfprdy = '1') then state := s4722;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4721; end if;
when s4722 => state := s4723; 	--15
	addfpsclr <= '0';
when s4723 => state := s4724; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4724 => 			--17
	if (addfprdy = '1') then state := s4725;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4724; end if;
when s4725 => state := s4726; 	--18
	addfpsclr <= '0';
when s4726 => state := s4727; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4727 => 			--20
	if (addfprdy = '1') then state := s4728;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4727; end if;
when s4728 => state := s4729; 	--21
	addfpsclr <= '0';
when s4729 => state := s4730; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (270, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4730 => state := s4731; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (478, 12)); -- offset LSB 430
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s4731 => state := s4732;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (479, 12)); -- offset MSB 431
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4732 => state := s4733; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4733 => 			--4
	if (fixed2floatrdy = '1') then state := s4734;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4733; end if;
when s4734 => state := s4735; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4735 => 			--6
	if (mulfprdy = '1') then state := s4736;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4735; end if;
when s4736 => state := s4737; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4737 => 			--8
	if (mulfprdy = '1') then state := s4738;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4737; end if;
when s4738 => state := s4739; 	--9
	mulfpsclr <= '0';
when s4739 => state := s4740; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4740 => 			--11
	if (mulfprdy = '1') then state := s4741;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4740; end if;
when s4741 => state := s4742; 	--12
	mulfpsclr <= '0';
when s4742 => state := s4743; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4743 => 			--14
	if (addfprdy = '1') then state := s4744;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4743; end if;
when s4744 => state := s4745; 	--15
	addfpsclr <= '0';
when s4745 => state := s4746; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4746 => 			--17
	if (addfprdy = '1') then state := s4747;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4746; end if;
when s4747 => state := s4748; 	--18
	addfpsclr <= '0';
when s4748 => state := s4749; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4749 => 			--20
	if (addfprdy = '1') then state := s4750;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4749; end if;
when s4750 => state := s4751; 	--21
	addfpsclr <= '0';
when s4751 => state := s4752; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (271, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4752 => state := s4753; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (480, 12)); -- offset LSB 432
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s4753 => state := s4754;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (481, 12)); -- offset MSB 433
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4754 => state := s4755; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4755 => 			--4
	if (fixed2floatrdy = '1') then state := s4756;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4755; end if;
when s4756 => state := s4757; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4757 => 			--6
	if (mulfprdy = '1') then state := s4758;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4757; end if;
when s4758 => state := s4759; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4759 => 			--8
	if (mulfprdy = '1') then state := s4760;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4759; end if;
when s4760 => state := s4761; 	--9
	mulfpsclr <= '0';
when s4761 => state := s4762; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4762 => 			--11
	if (mulfprdy = '1') then state := s4763;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4762; end if;
when s4763 => state := s4764; 	--12
	mulfpsclr <= '0';
when s4764 => state := s4765; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4765 => 			--14
	if (addfprdy = '1') then state := s4766;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4765; end if;
when s4766 => state := s4767; 	--15
	addfpsclr <= '0';
when s4767 => state := s4768; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4768 => 			--17
	if (addfprdy = '1') then state := s4769;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4768; end if;
when s4769 => state := s4770; 	--18
	addfpsclr <= '0';
when s4770 => state := s4771; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4771 => 			--20
	if (addfprdy = '1') then state := s4772;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4771; end if;
when s4772 => state := s4773; 	--21
	addfpsclr <= '0';
when s4773 => state := s4774; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (272, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4774 => state := s4775; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (482, 12)); -- offset LSB 434
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s4775 => state := s4776;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (483, 12)); -- offset MSB 435
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4776 => state := s4777; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4777 => 			--4
	if (fixed2floatrdy = '1') then state := s4778;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4777; end if;
when s4778 => state := s4779; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4779 => 			--6
	if (mulfprdy = '1') then state := s4780;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4779; end if;
when s4780 => state := s4781; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4781 => 			--8
	if (mulfprdy = '1') then state := s4782;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4781; end if;
when s4782 => state := s4783; 	--9
	mulfpsclr <= '0';
when s4783 => state := s4784; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4784 => 			--11
	if (mulfprdy = '1') then state := s4785;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4784; end if;
when s4785 => state := s4786; 	--12
	mulfpsclr <= '0';
when s4786 => state := s4787; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4787 => 			--14
	if (addfprdy = '1') then state := s4788;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4787; end if;
when s4788 => state := s4789; 	--15
	addfpsclr <= '0';
when s4789 => state := s4790; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4790 => 			--17
	if (addfprdy = '1') then state := s4791;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4790; end if;
when s4791 => state := s4792; 	--18
	addfpsclr <= '0';
when s4792 => state := s4793; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4793 => 			--20
	if (addfprdy = '1') then state := s4794;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4793; end if;
when s4794 => state := s4795; 	--21
	addfpsclr <= '0';
when s4795 => state := s4796; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (273, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4796 => state := s4797; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (484, 12)); -- offset LSB 436
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s4797 => state := s4798;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (485, 12)); -- offset MSB 437
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4798 => state := s4799; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4799 => 			--4
	if (fixed2floatrdy = '1') then state := s4800;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4799; end if;
when s4800 => state := s4801; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4801 => 			--6
	if (mulfprdy = '1') then state := s4802;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4801; end if;
when s4802 => state := s4803; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4803 => 			--8
	if (mulfprdy = '1') then state := s4804;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4803; end if;
when s4804 => state := s4805; 	--9
	mulfpsclr <= '0';
when s4805 => state := s4806; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4806 => 			--11
	if (mulfprdy = '1') then state := s4807;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4806; end if;
when s4807 => state := s4808; 	--12
	mulfpsclr <= '0';
when s4808 => state := s4809; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4809 => 			--14
	if (addfprdy = '1') then state := s4810;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4809; end if;
when s4810 => state := s4811; 	--15
	addfpsclr <= '0';
when s4811 => state := s4812; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4812 => 			--17
	if (addfprdy = '1') then state := s4813;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4812; end if;
when s4813 => state := s4814; 	--18
	addfpsclr <= '0';
when s4814 => state := s4815; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4815 => 			--20
	if (addfprdy = '1') then state := s4816;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4815; end if;
when s4816 => state := s4817; 	--21
	addfpsclr <= '0';
when s4817 => state := s4818; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (274, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4818 => state := s4819; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (486, 12)); -- offset LSB 438
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s4819 => state := s4820;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (487, 12)); -- offset MSB 439
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4820 => state := s4821; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4821 => 			--4
	if (fixed2floatrdy = '1') then state := s4822;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4821; end if;
when s4822 => state := s4823; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4823 => 			--6
	if (mulfprdy = '1') then state := s4824;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4823; end if;
when s4824 => state := s4825; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4825 => 			--8
	if (mulfprdy = '1') then state := s4826;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4825; end if;
when s4826 => state := s4827; 	--9
	mulfpsclr <= '0';
when s4827 => state := s4828; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4828 => 			--11
	if (mulfprdy = '1') then state := s4829;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4828; end if;
when s4829 => state := s4830; 	--12
	mulfpsclr <= '0';
when s4830 => state := s4831; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4831 => 			--14
	if (addfprdy = '1') then state := s4832;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4831; end if;
when s4832 => state := s4833; 	--15
	addfpsclr <= '0';
when s4833 => state := s4834; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4834 => 			--17
	if (addfprdy = '1') then state := s4835;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4834; end if;
when s4835 => state := s4836; 	--18
	addfpsclr <= '0';
when s4836 => state := s4837; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4837 => 			--20
	if (addfprdy = '1') then state := s4838;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4837; end if;
when s4838 => state := s4839; 	--21
	addfpsclr <= '0';
when s4839 => state := s4840; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (275, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4840 => state := s4841; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (488, 12)); -- offset LSB 440
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s4841 => state := s4842;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (489, 12)); -- offset MSB 441
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4842 => state := s4843; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4843 => 			--4
	if (fixed2floatrdy = '1') then state := s4844;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4843; end if;
when s4844 => state := s4845; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4845 => 			--6
	if (mulfprdy = '1') then state := s4846;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4845; end if;
when s4846 => state := s4847; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4847 => 			--8
	if (mulfprdy = '1') then state := s4848;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4847; end if;
when s4848 => state := s4849; 	--9
	mulfpsclr <= '0';
when s4849 => state := s4850; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4850 => 			--11
	if (mulfprdy = '1') then state := s4851;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4850; end if;
when s4851 => state := s4852; 	--12
	mulfpsclr <= '0';
when s4852 => state := s4853; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4853 => 			--14
	if (addfprdy = '1') then state := s4854;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4853; end if;
when s4854 => state := s4855; 	--15
	addfpsclr <= '0';
when s4855 => state := s4856; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4856 => 			--17
	if (addfprdy = '1') then state := s4857;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4856; end if;
when s4857 => state := s4858; 	--18
	addfpsclr <= '0';
when s4858 => state := s4859; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4859 => 			--20
	if (addfprdy = '1') then state := s4860;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4859; end if;
when s4860 => state := s4861; 	--21
	addfpsclr <= '0';
when s4861 => state := s4862; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (276, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4862 => state := s4863; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (490, 12)); -- offset LSB 442
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s4863 => state := s4864;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (491, 12)); -- offset MSB 443
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4864 => state := s4865; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4865 => 			--4
	if (fixed2floatrdy = '1') then state := s4866;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4865; end if;
when s4866 => state := s4867; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4867 => 			--6
	if (mulfprdy = '1') then state := s4868;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4867; end if;
when s4868 => state := s4869; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4869 => 			--8
	if (mulfprdy = '1') then state := s4870;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4869; end if;
when s4870 => state := s4871; 	--9
	mulfpsclr <= '0';
when s4871 => state := s4872; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4872 => 			--11
	if (mulfprdy = '1') then state := s4873;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4872; end if;
when s4873 => state := s4874; 	--12
	mulfpsclr <= '0';
when s4874 => state := s4875; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4875 => 			--14
	if (addfprdy = '1') then state := s4876;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4875; end if;
when s4876 => state := s4877; 	--15
	addfpsclr <= '0';
when s4877 => state := s4878; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4878 => 			--17
	if (addfprdy = '1') then state := s4879;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4878; end if;
when s4879 => state := s4880; 	--18
	addfpsclr <= '0';
when s4880 => state := s4881; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4881 => 			--20
	if (addfprdy = '1') then state := s4882;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4881; end if;
when s4882 => state := s4883; 	--21
	addfpsclr <= '0';
when s4883 => state := s4884; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (277, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4884 => state := s4885; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (492, 12)); -- offset LSB 444
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s4885 => state := s4886;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (493, 12)); -- offset MSB 445
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4886 => state := s4887; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4887 => 			--4
	if (fixed2floatrdy = '1') then state := s4888;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4887; end if;
when s4888 => state := s4889; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4889 => 			--6
	if (mulfprdy = '1') then state := s4890;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4889; end if;
when s4890 => state := s4891; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4891 => 			--8
	if (mulfprdy = '1') then state := s4892;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4891; end if;
when s4892 => state := s4893; 	--9
	mulfpsclr <= '0';
when s4893 => state := s4894; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4894 => 			--11
	if (mulfprdy = '1') then state := s4895;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4894; end if;
when s4895 => state := s4896; 	--12
	mulfpsclr <= '0';
when s4896 => state := s4897; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4897 => 			--14
	if (addfprdy = '1') then state := s4898;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4897; end if;
when s4898 => state := s4899; 	--15
	addfpsclr <= '0';
when s4899 => state := s4900; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4900 => 			--17
	if (addfprdy = '1') then state := s4901;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4900; end if;
when s4901 => state := s4902; 	--18
	addfpsclr <= '0';
when s4902 => state := s4903; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4903 => 			--20
	if (addfprdy = '1') then state := s4904;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4903; end if;
when s4904 => state := s4905; 	--21
	addfpsclr <= '0';
when s4905 => state := s4906; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (278, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4906 => state := s4907; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (494, 12)); -- offset LSB 446
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s4907 => state := s4908;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (495, 12)); -- offset MSB 447
	addra <= std_logic_vector (to_unsigned (6, 10)); -- OCCrowI 6
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4908 => state := s4909; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4909 => 			--4
	if (fixed2floatrdy = '1') then state := s4910;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4909; end if;
when s4910 => state := s4911; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4911 => 			--6
	if (mulfprdy = '1') then state := s4912;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4911; end if;
when s4912 => state := s4913; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4913 => 			--8
	if (mulfprdy = '1') then state := s4914;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4913; end if;
when s4914 => state := s4915; 	--9
	mulfpsclr <= '0';
when s4915 => state := s4916; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4916 => 			--11
	if (mulfprdy = '1') then state := s4917;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4916; end if;
when s4917 => state := s4918; 	--12
	mulfpsclr <= '0';
when s4918 => state := s4919; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4919 => 			--14
	if (addfprdy = '1') then state := s4920;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4919; end if;
when s4920 => state := s4921; 	--15
	addfpsclr <= '0';
when s4921 => state := s4922; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4922 => 			--17
	if (addfprdy = '1') then state := s4923;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4922; end if;
when s4923 => state := s4924; 	--18
	addfpsclr <= '0';
when s4924 => state := s4925; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4925 => 			--20
	if (addfprdy = '1') then state := s4926;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4925; end if;
when s4926 => state := s4927; 	--21
	addfpsclr <= '0';
when s4927 => state := s4928; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (279, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4928 => state := s4929; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (496, 12)); -- offset LSB 448
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s4929 => state := s4930;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (497, 12)); -- offset MSB 449
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4930 => state := s4931; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4931 => 			--4
	if (fixed2floatrdy = '1') then state := s4932;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4931; end if;
when s4932 => state := s4933; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4933 => 			--6
	if (mulfprdy = '1') then state := s4934;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4933; end if;
when s4934 => state := s4935; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4935 => 			--8
	if (mulfprdy = '1') then state := s4936;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4935; end if;
when s4936 => state := s4937; 	--9
	mulfpsclr <= '0';
when s4937 => state := s4938; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4938 => 			--11
	if (mulfprdy = '1') then state := s4939;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4938; end if;
when s4939 => state := s4940; 	--12
	mulfpsclr <= '0';
when s4940 => state := s4941; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4941 => 			--14
	if (addfprdy = '1') then state := s4942;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4941; end if;
when s4942 => state := s4943; 	--15
	addfpsclr <= '0';
when s4943 => state := s4944; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4944 => 			--17
	if (addfprdy = '1') then state := s4945;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4944; end if;
when s4945 => state := s4946; 	--18
	addfpsclr <= '0';
when s4946 => state := s4947; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4947 => 			--20
	if (addfprdy = '1') then state := s4948;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4947; end if;
when s4948 => state := s4949; 	--21
	addfpsclr <= '0';
when s4949 => state := s4950; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (280, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4950 => state := s4951; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (498, 12)); -- offset LSB 450
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s4951 => state := s4952;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (499, 12)); -- offset MSB 451
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4952 => state := s4953; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4953 => 			--4
	if (fixed2floatrdy = '1') then state := s4954;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4953; end if;
when s4954 => state := s4955; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4955 => 			--6
	if (mulfprdy = '1') then state := s4956;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4955; end if;
when s4956 => state := s4957; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4957 => 			--8
	if (mulfprdy = '1') then state := s4958;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4957; end if;
when s4958 => state := s4959; 	--9
	mulfpsclr <= '0';
when s4959 => state := s4960; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4960 => 			--11
	if (mulfprdy = '1') then state := s4961;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4960; end if;
when s4961 => state := s4962; 	--12
	mulfpsclr <= '0';
when s4962 => state := s4963; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4963 => 			--14
	if (addfprdy = '1') then state := s4964;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4963; end if;
when s4964 => state := s4965; 	--15
	addfpsclr <= '0';
when s4965 => state := s4966; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4966 => 			--17
	if (addfprdy = '1') then state := s4967;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4966; end if;
when s4967 => state := s4968; 	--18
	addfpsclr <= '0';
when s4968 => state := s4969; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4969 => 			--20
	if (addfprdy = '1') then state := s4970;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4969; end if;
when s4970 => state := s4971; 	--21
	addfpsclr <= '0';
when s4971 => state := s4972; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (281, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4972 => state := s4973; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (500, 12)); -- offset LSB 452
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s4973 => state := s4974;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (501, 12)); -- offset MSB 453
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4974 => state := s4975; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4975 => 			--4
	if (fixed2floatrdy = '1') then state := s4976;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4975; end if;
when s4976 => state := s4977; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4977 => 			--6
	if (mulfprdy = '1') then state := s4978;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4977; end if;
when s4978 => state := s4979; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s4979 => 			--8
	if (mulfprdy = '1') then state := s4980;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4979; end if;
when s4980 => state := s4981; 	--9
	mulfpsclr <= '0';
when s4981 => state := s4982; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s4982 => 			--11
	if (mulfprdy = '1') then state := s4983;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4982; end if;
when s4983 => state := s4984; 	--12
	mulfpsclr <= '0';
when s4984 => state := s4985; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s4985 => 			--14
	if (addfprdy = '1') then state := s4986;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4985; end if;
when s4986 => state := s4987; 	--15
	addfpsclr <= '0';
when s4987 => state := s4988; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s4988 => 			--17
	if (addfprdy = '1') then state := s4989;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4988; end if;
when s4989 => state := s4990; 	--18
	addfpsclr <= '0';
when s4990 => state := s4991; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s4991 => 			--20
	if (addfprdy = '1') then state := s4992;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s4991; end if;
when s4992 => state := s4993; 	--21
	addfpsclr <= '0';
when s4993 => state := s4994; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (282, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s4994 => state := s4995; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (502, 12)); -- offset LSB 454
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s4995 => state := s4996;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (503, 12)); -- offset MSB 455
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s4996 => state := s4997; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s4997 => 			--4
	if (fixed2floatrdy = '1') then state := s4998;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s4997; end if;
when s4998 => state := s4999; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s4999 => 			--6
	if (mulfprdy = '1') then state := s5000;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s4999; end if;
when s5000 => state := s5001; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5001 => 			--8
	if (mulfprdy = '1') then state := s5002;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5001; end if;
when s5002 => state := s5003; 	--9
	mulfpsclr <= '0';
when s5003 => state := s5004; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5004 => 			--11
	if (mulfprdy = '1') then state := s5005;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5004; end if;
when s5005 => state := s5006; 	--12
	mulfpsclr <= '0';
when s5006 => state := s5007; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5007 => 			--14
	if (addfprdy = '1') then state := s5008;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5007; end if;
when s5008 => state := s5009; 	--15
	addfpsclr <= '0';
when s5009 => state := s5010; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5010 => 			--17
	if (addfprdy = '1') then state := s5011;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5010; end if;
when s5011 => state := s5012; 	--18
	addfpsclr <= '0';
when s5012 => state := s5013; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5013 => 			--20
	if (addfprdy = '1') then state := s5014;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5013; end if;
when s5014 => state := s5015; 	--21
	addfpsclr <= '0';
when s5015 => state := s5016; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (283, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5016 => state := s5017; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (504, 12)); -- offset LSB 456
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s5017 => state := s5018;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (505, 12)); -- offset MSB 457
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5018 => state := s5019; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5019 => 			--4
	if (fixed2floatrdy = '1') then state := s5020;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5019; end if;
when s5020 => state := s5021; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5021 => 			--6
	if (mulfprdy = '1') then state := s5022;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5021; end if;
when s5022 => state := s5023; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5023 => 			--8
	if (mulfprdy = '1') then state := s5024;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5023; end if;
when s5024 => state := s5025; 	--9
	mulfpsclr <= '0';
when s5025 => state := s5026; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5026 => 			--11
	if (mulfprdy = '1') then state := s5027;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5026; end if;
when s5027 => state := s5028; 	--12
	mulfpsclr <= '0';
when s5028 => state := s5029; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5029 => 			--14
	if (addfprdy = '1') then state := s5030;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5029; end if;
when s5030 => state := s5031; 	--15
	addfpsclr <= '0';
when s5031 => state := s5032; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5032 => 			--17
	if (addfprdy = '1') then state := s5033;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5032; end if;
when s5033 => state := s5034; 	--18
	addfpsclr <= '0';
when s5034 => state := s5035; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5035 => 			--20
	if (addfprdy = '1') then state := s5036;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5035; end if;
when s5036 => state := s5037; 	--21
	addfpsclr <= '0';
when s5037 => state := s5038; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (284, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5038 => state := s5039; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (506, 12)); -- offset LSB 458
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s5039 => state := s5040;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (507, 12)); -- offset MSB 459
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5040 => state := s5041; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5041 => 			--4
	if (fixed2floatrdy = '1') then state := s5042;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5041; end if;
when s5042 => state := s5043; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5043 => 			--6
	if (mulfprdy = '1') then state := s5044;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5043; end if;
when s5044 => state := s5045; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5045 => 			--8
	if (mulfprdy = '1') then state := s5046;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5045; end if;
when s5046 => state := s5047; 	--9
	mulfpsclr <= '0';
when s5047 => state := s5048; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5048 => 			--11
	if (mulfprdy = '1') then state := s5049;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5048; end if;
when s5049 => state := s5050; 	--12
	mulfpsclr <= '0';
when s5050 => state := s5051; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5051 => 			--14
	if (addfprdy = '1') then state := s5052;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5051; end if;
when s5052 => state := s5053; 	--15
	addfpsclr <= '0';
when s5053 => state := s5054; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5054 => 			--17
	if (addfprdy = '1') then state := s5055;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5054; end if;
when s5055 => state := s5056; 	--18
	addfpsclr <= '0';
when s5056 => state := s5057; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5057 => 			--20
	if (addfprdy = '1') then state := s5058;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5057; end if;
when s5058 => state := s5059; 	--21
	addfpsclr <= '0';
when s5059 => state := s5060; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (285, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5060 => state := s5061; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (508, 12)); -- offset LSB 460
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s5061 => state := s5062;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (509, 12)); -- offset MSB 461
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5062 => state := s5063; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5063 => 			--4
	if (fixed2floatrdy = '1') then state := s5064;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5063; end if;
when s5064 => state := s5065; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5065 => 			--6
	if (mulfprdy = '1') then state := s5066;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5065; end if;
when s5066 => state := s5067; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5067 => 			--8
	if (mulfprdy = '1') then state := s5068;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5067; end if;
when s5068 => state := s5069; 	--9
	mulfpsclr <= '0';
when s5069 => state := s5070; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5070 => 			--11
	if (mulfprdy = '1') then state := s5071;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5070; end if;
when s5071 => state := s5072; 	--12
	mulfpsclr <= '0';
when s5072 => state := s5073; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5073 => 			--14
	if (addfprdy = '1') then state := s5074;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5073; end if;
when s5074 => state := s5075; 	--15
	addfpsclr <= '0';
when s5075 => state := s5076; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5076 => 			--17
	if (addfprdy = '1') then state := s5077;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5076; end if;
when s5077 => state := s5078; 	--18
	addfpsclr <= '0';
when s5078 => state := s5079; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5079 => 			--20
	if (addfprdy = '1') then state := s5080;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5079; end if;
when s5080 => state := s5081; 	--21
	addfpsclr <= '0';
when s5081 => state := s5082; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (286, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5082 => state := s5083; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (510, 12)); -- offset LSB 462
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s5083 => state := s5084;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (511, 12)); -- offset MSB 463
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5084 => state := s5085; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5085 => 			--4
	if (fixed2floatrdy = '1') then state := s5086;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5085; end if;
when s5086 => state := s5087; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5087 => 			--6
	if (mulfprdy = '1') then state := s5088;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5087; end if;
when s5088 => state := s5089; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5089 => 			--8
	if (mulfprdy = '1') then state := s5090;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5089; end if;
when s5090 => state := s5091; 	--9
	mulfpsclr <= '0';
when s5091 => state := s5092; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5092 => 			--11
	if (mulfprdy = '1') then state := s5093;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5092; end if;
when s5093 => state := s5094; 	--12
	mulfpsclr <= '0';
when s5094 => state := s5095; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5095 => 			--14
	if (addfprdy = '1') then state := s5096;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5095; end if;
when s5096 => state := s5097; 	--15
	addfpsclr <= '0';
when s5097 => state := s5098; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5098 => 			--17
	if (addfprdy = '1') then state := s5099;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5098; end if;
when s5099 => state := s5100; 	--18
	addfpsclr <= '0';
when s5100 => state := s5101; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5101 => 			--20
	if (addfprdy = '1') then state := s5102;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5101; end if;
when s5102 => state := s5103; 	--21
	addfpsclr <= '0';
when s5103 => state := s5104; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (287, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5104 => state := s5105; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (512, 12)); -- offset LSB 464
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s5105 => state := s5106;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (513, 12)); -- offset MSB 465
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5106 => state := s5107; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5107 => 			--4
	if (fixed2floatrdy = '1') then state := s5108;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5107; end if;
when s5108 => state := s5109; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5109 => 			--6
	if (mulfprdy = '1') then state := s5110;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5109; end if;
when s5110 => state := s5111; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5111 => 			--8
	if (mulfprdy = '1') then state := s5112;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5111; end if;
when s5112 => state := s5113; 	--9
	mulfpsclr <= '0';
when s5113 => state := s5114; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5114 => 			--11
	if (mulfprdy = '1') then state := s5115;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5114; end if;
when s5115 => state := s5116; 	--12
	mulfpsclr <= '0';
when s5116 => state := s5117; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5117 => 			--14
	if (addfprdy = '1') then state := s5118;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5117; end if;
when s5118 => state := s5119; 	--15
	addfpsclr <= '0';
when s5119 => state := s5120; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5120 => 			--17
	if (addfprdy = '1') then state := s5121;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5120; end if;
when s5121 => state := s5122; 	--18
	addfpsclr <= '0';
when s5122 => state := s5123; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5123 => 			--20
	if (addfprdy = '1') then state := s5124;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5123; end if;
when s5124 => state := s5125; 	--21
	addfpsclr <= '0';
when s5125 => state := s5126; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (288, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5126 => state := s5127; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (514, 12)); -- offset LSB 466
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s5127 => state := s5128;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (515, 12)); -- offset MSB 467
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5128 => state := s5129; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5129 => 			--4
	if (fixed2floatrdy = '1') then state := s5130;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5129; end if;
when s5130 => state := s5131; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5131 => 			--6
	if (mulfprdy = '1') then state := s5132;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5131; end if;
when s5132 => state := s5133; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5133 => 			--8
	if (mulfprdy = '1') then state := s5134;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5133; end if;
when s5134 => state := s5135; 	--9
	mulfpsclr <= '0';
when s5135 => state := s5136; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5136 => 			--11
	if (mulfprdy = '1') then state := s5137;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5136; end if;
when s5137 => state := s5138; 	--12
	mulfpsclr <= '0';
when s5138 => state := s5139; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5139 => 			--14
	if (addfprdy = '1') then state := s5140;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5139; end if;
when s5140 => state := s5141; 	--15
	addfpsclr <= '0';
when s5141 => state := s5142; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5142 => 			--17
	if (addfprdy = '1') then state := s5143;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5142; end if;
when s5143 => state := s5144; 	--18
	addfpsclr <= '0';
when s5144 => state := s5145; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5145 => 			--20
	if (addfprdy = '1') then state := s5146;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5145; end if;
when s5146 => state := s5147; 	--21
	addfpsclr <= '0';
when s5147 => state := s5148; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (289, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5148 => state := s5149; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (516, 12)); -- offset LSB 468
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s5149 => state := s5150;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (517, 12)); -- offset MSB 469
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5150 => state := s5151; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5151 => 			--4
	if (fixed2floatrdy = '1') then state := s5152;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5151; end if;
when s5152 => state := s5153; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5153 => 			--6
	if (mulfprdy = '1') then state := s5154;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5153; end if;
when s5154 => state := s5155; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5155 => 			--8
	if (mulfprdy = '1') then state := s5156;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5155; end if;
when s5156 => state := s5157; 	--9
	mulfpsclr <= '0';
when s5157 => state := s5158; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5158 => 			--11
	if (mulfprdy = '1') then state := s5159;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5158; end if;
when s5159 => state := s5160; 	--12
	mulfpsclr <= '0';
when s5160 => state := s5161; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5161 => 			--14
	if (addfprdy = '1') then state := s5162;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5161; end if;
when s5162 => state := s5163; 	--15
	addfpsclr <= '0';
when s5163 => state := s5164; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5164 => 			--17
	if (addfprdy = '1') then state := s5165;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5164; end if;
when s5165 => state := s5166; 	--18
	addfpsclr <= '0';
when s5166 => state := s5167; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5167 => 			--20
	if (addfprdy = '1') then state := s5168;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5167; end if;
when s5168 => state := s5169; 	--21
	addfpsclr <= '0';
when s5169 => state := s5170; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (290, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5170 => state := s5171; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (518, 12)); -- offset LSB 470
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s5171 => state := s5172;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (519, 12)); -- offset MSB 471
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5172 => state := s5173; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5173 => 			--4
	if (fixed2floatrdy = '1') then state := s5174;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5173; end if;
when s5174 => state := s5175; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5175 => 			--6
	if (mulfprdy = '1') then state := s5176;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5175; end if;
when s5176 => state := s5177; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5177 => 			--8
	if (mulfprdy = '1') then state := s5178;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5177; end if;
when s5178 => state := s5179; 	--9
	mulfpsclr <= '0';
when s5179 => state := s5180; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5180 => 			--11
	if (mulfprdy = '1') then state := s5181;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5180; end if;
when s5181 => state := s5182; 	--12
	mulfpsclr <= '0';
when s5182 => state := s5183; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5183 => 			--14
	if (addfprdy = '1') then state := s5184;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5183; end if;
when s5184 => state := s5185; 	--15
	addfpsclr <= '0';
when s5185 => state := s5186; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5186 => 			--17
	if (addfprdy = '1') then state := s5187;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5186; end if;
when s5187 => state := s5188; 	--18
	addfpsclr <= '0';
when s5188 => state := s5189; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5189 => 			--20
	if (addfprdy = '1') then state := s5190;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5189; end if;
when s5190 => state := s5191; 	--21
	addfpsclr <= '0';
when s5191 => state := s5192; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (291, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5192 => state := s5193; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (520, 12)); -- offset LSB 472
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s5193 => state := s5194;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (521, 12)); -- offset MSB 473
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5194 => state := s5195; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5195 => 			--4
	if (fixed2floatrdy = '1') then state := s5196;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5195; end if;
when s5196 => state := s5197; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5197 => 			--6
	if (mulfprdy = '1') then state := s5198;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5197; end if;
when s5198 => state := s5199; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5199 => 			--8
	if (mulfprdy = '1') then state := s5200;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5199; end if;
when s5200 => state := s5201; 	--9
	mulfpsclr <= '0';
when s5201 => state := s5202; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5202 => 			--11
	if (mulfprdy = '1') then state := s5203;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5202; end if;
when s5203 => state := s5204; 	--12
	mulfpsclr <= '0';
when s5204 => state := s5205; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5205 => 			--14
	if (addfprdy = '1') then state := s5206;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5205; end if;
when s5206 => state := s5207; 	--15
	addfpsclr <= '0';
when s5207 => state := s5208; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5208 => 			--17
	if (addfprdy = '1') then state := s5209;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5208; end if;
when s5209 => state := s5210; 	--18
	addfpsclr <= '0';
when s5210 => state := s5211; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5211 => 			--20
	if (addfprdy = '1') then state := s5212;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5211; end if;
when s5212 => state := s5213; 	--21
	addfpsclr <= '0';
when s5213 => state := s5214; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (292, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5214 => state := s5215; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (522, 12)); -- offset LSB 474
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s5215 => state := s5216;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (523, 12)); -- offset MSB 475
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5216 => state := s5217; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5217 => 			--4
	if (fixed2floatrdy = '1') then state := s5218;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5217; end if;
when s5218 => state := s5219; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5219 => 			--6
	if (mulfprdy = '1') then state := s5220;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5219; end if;
when s5220 => state := s5221; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5221 => 			--8
	if (mulfprdy = '1') then state := s5222;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5221; end if;
when s5222 => state := s5223; 	--9
	mulfpsclr <= '0';
when s5223 => state := s5224; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5224 => 			--11
	if (mulfprdy = '1') then state := s5225;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5224; end if;
when s5225 => state := s5226; 	--12
	mulfpsclr <= '0';
when s5226 => state := s5227; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5227 => 			--14
	if (addfprdy = '1') then state := s5228;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5227; end if;
when s5228 => state := s5229; 	--15
	addfpsclr <= '0';
when s5229 => state := s5230; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5230 => 			--17
	if (addfprdy = '1') then state := s5231;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5230; end if;
when s5231 => state := s5232; 	--18
	addfpsclr <= '0';
when s5232 => state := s5233; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5233 => 			--20
	if (addfprdy = '1') then state := s5234;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5233; end if;
when s5234 => state := s5235; 	--21
	addfpsclr <= '0';
when s5235 => state := s5236; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (293, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5236 => state := s5237; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (524, 12)); -- offset LSB 476
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s5237 => state := s5238;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (525, 12)); -- offset MSB 477
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5238 => state := s5239; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5239 => 			--4
	if (fixed2floatrdy = '1') then state := s5240;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5239; end if;
when s5240 => state := s5241; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5241 => 			--6
	if (mulfprdy = '1') then state := s5242;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5241; end if;
when s5242 => state := s5243; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5243 => 			--8
	if (mulfprdy = '1') then state := s5244;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5243; end if;
when s5244 => state := s5245; 	--9
	mulfpsclr <= '0';
when s5245 => state := s5246; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5246 => 			--11
	if (mulfprdy = '1') then state := s5247;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5246; end if;
when s5247 => state := s5248; 	--12
	mulfpsclr <= '0';
when s5248 => state := s5249; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5249 => 			--14
	if (addfprdy = '1') then state := s5250;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5249; end if;
when s5250 => state := s5251; 	--15
	addfpsclr <= '0';
when s5251 => state := s5252; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5252 => 			--17
	if (addfprdy = '1') then state := s5253;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5252; end if;
when s5253 => state := s5254; 	--18
	addfpsclr <= '0';
when s5254 => state := s5255; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5255 => 			--20
	if (addfprdy = '1') then state := s5256;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5255; end if;
when s5256 => state := s5257; 	--21
	addfpsclr <= '0';
when s5257 => state := s5258; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (294, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5258 => state := s5259; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (526, 12)); -- offset LSB 478
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s5259 => state := s5260;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (527, 12)); -- offset MSB 479
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5260 => state := s5261; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5261 => 			--4
	if (fixed2floatrdy = '1') then state := s5262;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5261; end if;
when s5262 => state := s5263; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5263 => 			--6
	if (mulfprdy = '1') then state := s5264;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5263; end if;
when s5264 => state := s5265; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5265 => 			--8
	if (mulfprdy = '1') then state := s5266;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5265; end if;
when s5266 => state := s5267; 	--9
	mulfpsclr <= '0';
when s5267 => state := s5268; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5268 => 			--11
	if (mulfprdy = '1') then state := s5269;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5268; end if;
when s5269 => state := s5270; 	--12
	mulfpsclr <= '0';
when s5270 => state := s5271; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5271 => 			--14
	if (addfprdy = '1') then state := s5272;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5271; end if;
when s5272 => state := s5273; 	--15
	addfpsclr <= '0';
when s5273 => state := s5274; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5274 => 			--17
	if (addfprdy = '1') then state := s5275;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5274; end if;
when s5275 => state := s5276; 	--18
	addfpsclr <= '0';
when s5276 => state := s5277; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5277 => 			--20
	if (addfprdy = '1') then state := s5278;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5277; end if;
when s5278 => state := s5279; 	--21
	addfpsclr <= '0';
when s5279 => state := s5280; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (295, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5280 => state := s5281; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (528, 12)); -- offset LSB 480
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s5281 => state := s5282;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (529, 12)); -- offset MSB 481
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5282 => state := s5283; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5283 => 			--4
	if (fixed2floatrdy = '1') then state := s5284;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5283; end if;
when s5284 => state := s5285; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5285 => 			--6
	if (mulfprdy = '1') then state := s5286;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5285; end if;
when s5286 => state := s5287; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5287 => 			--8
	if (mulfprdy = '1') then state := s5288;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5287; end if;
when s5288 => state := s5289; 	--9
	mulfpsclr <= '0';
when s5289 => state := s5290; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5290 => 			--11
	if (mulfprdy = '1') then state := s5291;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5290; end if;
when s5291 => state := s5292; 	--12
	mulfpsclr <= '0';
when s5292 => state := s5293; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5293 => 			--14
	if (addfprdy = '1') then state := s5294;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5293; end if;
when s5294 => state := s5295; 	--15
	addfpsclr <= '0';
when s5295 => state := s5296; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5296 => 			--17
	if (addfprdy = '1') then state := s5297;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5296; end if;
when s5297 => state := s5298; 	--18
	addfpsclr <= '0';
when s5298 => state := s5299; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5299 => 			--20
	if (addfprdy = '1') then state := s5300;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5299; end if;
when s5300 => state := s5301; 	--21
	addfpsclr <= '0';
when s5301 => state := s5302; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (296, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5302 => state := s5303; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (530, 12)); -- offset LSB 482
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s5303 => state := s5304;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (531, 12)); -- offset MSB 483
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5304 => state := s5305; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5305 => 			--4
	if (fixed2floatrdy = '1') then state := s5306;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5305; end if;
when s5306 => state := s5307; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5307 => 			--6
	if (mulfprdy = '1') then state := s5308;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5307; end if;
when s5308 => state := s5309; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5309 => 			--8
	if (mulfprdy = '1') then state := s5310;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5309; end if;
when s5310 => state := s5311; 	--9
	mulfpsclr <= '0';
when s5311 => state := s5312; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5312 => 			--11
	if (mulfprdy = '1') then state := s5313;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5312; end if;
when s5313 => state := s5314; 	--12
	mulfpsclr <= '0';
when s5314 => state := s5315; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5315 => 			--14
	if (addfprdy = '1') then state := s5316;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5315; end if;
when s5316 => state := s5317; 	--15
	addfpsclr <= '0';
when s5317 => state := s5318; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5318 => 			--17
	if (addfprdy = '1') then state := s5319;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5318; end if;
when s5319 => state := s5320; 	--18
	addfpsclr <= '0';
when s5320 => state := s5321; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5321 => 			--20
	if (addfprdy = '1') then state := s5322;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5321; end if;
when s5322 => state := s5323; 	--21
	addfpsclr <= '0';
when s5323 => state := s5324; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (297, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5324 => state := s5325; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (532, 12)); -- offset LSB 484
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s5325 => state := s5326;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (533, 12)); -- offset MSB 485
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5326 => state := s5327; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5327 => 			--4
	if (fixed2floatrdy = '1') then state := s5328;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5327; end if;
when s5328 => state := s5329; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5329 => 			--6
	if (mulfprdy = '1') then state := s5330;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5329; end if;
when s5330 => state := s5331; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5331 => 			--8
	if (mulfprdy = '1') then state := s5332;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5331; end if;
when s5332 => state := s5333; 	--9
	mulfpsclr <= '0';
when s5333 => state := s5334; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5334 => 			--11
	if (mulfprdy = '1') then state := s5335;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5334; end if;
when s5335 => state := s5336; 	--12
	mulfpsclr <= '0';
when s5336 => state := s5337; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5337 => 			--14
	if (addfprdy = '1') then state := s5338;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5337; end if;
when s5338 => state := s5339; 	--15
	addfpsclr <= '0';
when s5339 => state := s5340; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5340 => 			--17
	if (addfprdy = '1') then state := s5341;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5340; end if;
when s5341 => state := s5342; 	--18
	addfpsclr <= '0';
when s5342 => state := s5343; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5343 => 			--20
	if (addfprdy = '1') then state := s5344;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5343; end if;
when s5344 => state := s5345; 	--21
	addfpsclr <= '0';
when s5345 => state := s5346; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (298, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5346 => state := s5347; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (534, 12)); -- offset LSB 486
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s5347 => state := s5348;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (535, 12)); -- offset MSB 487
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5348 => state := s5349; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5349 => 			--4
	if (fixed2floatrdy = '1') then state := s5350;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5349; end if;
when s5350 => state := s5351; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5351 => 			--6
	if (mulfprdy = '1') then state := s5352;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5351; end if;
when s5352 => state := s5353; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5353 => 			--8
	if (mulfprdy = '1') then state := s5354;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5353; end if;
when s5354 => state := s5355; 	--9
	mulfpsclr <= '0';
when s5355 => state := s5356; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5356 => 			--11
	if (mulfprdy = '1') then state := s5357;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5356; end if;
when s5357 => state := s5358; 	--12
	mulfpsclr <= '0';
when s5358 => state := s5359; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5359 => 			--14
	if (addfprdy = '1') then state := s5360;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5359; end if;
when s5360 => state := s5361; 	--15
	addfpsclr <= '0';
when s5361 => state := s5362; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5362 => 			--17
	if (addfprdy = '1') then state := s5363;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5362; end if;
when s5363 => state := s5364; 	--18
	addfpsclr <= '0';
when s5364 => state := s5365; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5365 => 			--20
	if (addfprdy = '1') then state := s5366;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5365; end if;
when s5366 => state := s5367; 	--21
	addfpsclr <= '0';
when s5367 => state := s5368; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (299, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5368 => state := s5369; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (536, 12)); -- offset LSB 488
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s5369 => state := s5370;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (537, 12)); -- offset MSB 489
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5370 => state := s5371; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5371 => 			--4
	if (fixed2floatrdy = '1') then state := s5372;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5371; end if;
when s5372 => state := s5373; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5373 => 			--6
	if (mulfprdy = '1') then state := s5374;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5373; end if;
when s5374 => state := s5375; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5375 => 			--8
	if (mulfprdy = '1') then state := s5376;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5375; end if;
when s5376 => state := s5377; 	--9
	mulfpsclr <= '0';
when s5377 => state := s5378; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5378 => 			--11
	if (mulfprdy = '1') then state := s5379;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5378; end if;
when s5379 => state := s5380; 	--12
	mulfpsclr <= '0';
when s5380 => state := s5381; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5381 => 			--14
	if (addfprdy = '1') then state := s5382;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5381; end if;
when s5382 => state := s5383; 	--15
	addfpsclr <= '0';
when s5383 => state := s5384; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5384 => 			--17
	if (addfprdy = '1') then state := s5385;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5384; end if;
when s5385 => state := s5386; 	--18
	addfpsclr <= '0';
when s5386 => state := s5387; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5387 => 			--20
	if (addfprdy = '1') then state := s5388;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5387; end if;
when s5388 => state := s5389; 	--21
	addfpsclr <= '0';
when s5389 => state := s5390; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (300, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5390 => state := s5391; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (538, 12)); -- offset LSB 490
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s5391 => state := s5392;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (539, 12)); -- offset MSB 491
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5392 => state := s5393; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5393 => 			--4
	if (fixed2floatrdy = '1') then state := s5394;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5393; end if;
when s5394 => state := s5395; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5395 => 			--6
	if (mulfprdy = '1') then state := s5396;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5395; end if;
when s5396 => state := s5397; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5397 => 			--8
	if (mulfprdy = '1') then state := s5398;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5397; end if;
when s5398 => state := s5399; 	--9
	mulfpsclr <= '0';
when s5399 => state := s5400; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5400 => 			--11
	if (mulfprdy = '1') then state := s5401;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5400; end if;
when s5401 => state := s5402; 	--12
	mulfpsclr <= '0';
when s5402 => state := s5403; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5403 => 			--14
	if (addfprdy = '1') then state := s5404;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5403; end if;
when s5404 => state := s5405; 	--15
	addfpsclr <= '0';
when s5405 => state := s5406; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5406 => 			--17
	if (addfprdy = '1') then state := s5407;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5406; end if;
when s5407 => state := s5408; 	--18
	addfpsclr <= '0';
when s5408 => state := s5409; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5409 => 			--20
	if (addfprdy = '1') then state := s5410;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5409; end if;
when s5410 => state := s5411; 	--21
	addfpsclr <= '0';
when s5411 => state := s5412; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (301, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5412 => state := s5413; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (540, 12)); -- offset LSB 492
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s5413 => state := s5414;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (541, 12)); -- offset MSB 493
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5414 => state := s5415; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5415 => 			--4
	if (fixed2floatrdy = '1') then state := s5416;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5415; end if;
when s5416 => state := s5417; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5417 => 			--6
	if (mulfprdy = '1') then state := s5418;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5417; end if;
when s5418 => state := s5419; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5419 => 			--8
	if (mulfprdy = '1') then state := s5420;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5419; end if;
when s5420 => state := s5421; 	--9
	mulfpsclr <= '0';
when s5421 => state := s5422; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5422 => 			--11
	if (mulfprdy = '1') then state := s5423;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5422; end if;
when s5423 => state := s5424; 	--12
	mulfpsclr <= '0';
when s5424 => state := s5425; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5425 => 			--14
	if (addfprdy = '1') then state := s5426;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5425; end if;
when s5426 => state := s5427; 	--15
	addfpsclr <= '0';
when s5427 => state := s5428; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5428 => 			--17
	if (addfprdy = '1') then state := s5429;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5428; end if;
when s5429 => state := s5430; 	--18
	addfpsclr <= '0';
when s5430 => state := s5431; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5431 => 			--20
	if (addfprdy = '1') then state := s5432;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5431; end if;
when s5432 => state := s5433; 	--21
	addfpsclr <= '0';
when s5433 => state := s5434; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (302, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5434 => state := s5435; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (542, 12)); -- offset LSB 494
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s5435 => state := s5436;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (543, 12)); -- offset MSB 495
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5436 => state := s5437; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5437 => 			--4
	if (fixed2floatrdy = '1') then state := s5438;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5437; end if;
when s5438 => state := s5439; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5439 => 			--6
	if (mulfprdy = '1') then state := s5440;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5439; end if;
when s5440 => state := s5441; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5441 => 			--8
	if (mulfprdy = '1') then state := s5442;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5441; end if;
when s5442 => state := s5443; 	--9
	mulfpsclr <= '0';
when s5443 => state := s5444; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5444 => 			--11
	if (mulfprdy = '1') then state := s5445;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5444; end if;
when s5445 => state := s5446; 	--12
	mulfpsclr <= '0';
when s5446 => state := s5447; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5447 => 			--14
	if (addfprdy = '1') then state := s5448;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5447; end if;
when s5448 => state := s5449; 	--15
	addfpsclr <= '0';
when s5449 => state := s5450; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5450 => 			--17
	if (addfprdy = '1') then state := s5451;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5450; end if;
when s5451 => state := s5452; 	--18
	addfpsclr <= '0';
when s5452 => state := s5453; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5453 => 			--20
	if (addfprdy = '1') then state := s5454;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5453; end if;
when s5454 => state := s5455; 	--21
	addfpsclr <= '0';
when s5455 => state := s5456; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (303, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5456 => state := s5457; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (544, 12)); -- offset LSB 496
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s5457 => state := s5458;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (545, 12)); -- offset MSB 497
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5458 => state := s5459; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5459 => 			--4
	if (fixed2floatrdy = '1') then state := s5460;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5459; end if;
when s5460 => state := s5461; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5461 => 			--6
	if (mulfprdy = '1') then state := s5462;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5461; end if;
when s5462 => state := s5463; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5463 => 			--8
	if (mulfprdy = '1') then state := s5464;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5463; end if;
when s5464 => state := s5465; 	--9
	mulfpsclr <= '0';
when s5465 => state := s5466; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5466 => 			--11
	if (mulfprdy = '1') then state := s5467;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5466; end if;
when s5467 => state := s5468; 	--12
	mulfpsclr <= '0';
when s5468 => state := s5469; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5469 => 			--14
	if (addfprdy = '1') then state := s5470;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5469; end if;
when s5470 => state := s5471; 	--15
	addfpsclr <= '0';
when s5471 => state := s5472; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5472 => 			--17
	if (addfprdy = '1') then state := s5473;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5472; end if;
when s5473 => state := s5474; 	--18
	addfpsclr <= '0';
when s5474 => state := s5475; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5475 => 			--20
	if (addfprdy = '1') then state := s5476;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5475; end if;
when s5476 => state := s5477; 	--21
	addfpsclr <= '0';
when s5477 => state := s5478; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (304, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5478 => state := s5479; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (546, 12)); -- offset LSB 498
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s5479 => state := s5480;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (547, 12)); -- offset MSB 499
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5480 => state := s5481; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5481 => 			--4
	if (fixed2floatrdy = '1') then state := s5482;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5481; end if;
when s5482 => state := s5483; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5483 => 			--6
	if (mulfprdy = '1') then state := s5484;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5483; end if;
when s5484 => state := s5485; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5485 => 			--8
	if (mulfprdy = '1') then state := s5486;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5485; end if;
when s5486 => state := s5487; 	--9
	mulfpsclr <= '0';
when s5487 => state := s5488; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5488 => 			--11
	if (mulfprdy = '1') then state := s5489;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5488; end if;
when s5489 => state := s5490; 	--12
	mulfpsclr <= '0';
when s5490 => state := s5491; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5491 => 			--14
	if (addfprdy = '1') then state := s5492;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5491; end if;
when s5492 => state := s5493; 	--15
	addfpsclr <= '0';
when s5493 => state := s5494; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5494 => 			--17
	if (addfprdy = '1') then state := s5495;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5494; end if;
when s5495 => state := s5496; 	--18
	addfpsclr <= '0';
when s5496 => state := s5497; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5497 => 			--20
	if (addfprdy = '1') then state := s5498;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5497; end if;
when s5498 => state := s5499; 	--21
	addfpsclr <= '0';
when s5499 => state := s5500; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (305, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5500 => state := s5501; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (548, 12)); -- offset LSB 500
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s5501 => state := s5502;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (549, 12)); -- offset MSB 501
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5502 => state := s5503; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5503 => 			--4
	if (fixed2floatrdy = '1') then state := s5504;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5503; end if;
when s5504 => state := s5505; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5505 => 			--6
	if (mulfprdy = '1') then state := s5506;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5505; end if;
when s5506 => state := s5507; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5507 => 			--8
	if (mulfprdy = '1') then state := s5508;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5507; end if;
when s5508 => state := s5509; 	--9
	mulfpsclr <= '0';
when s5509 => state := s5510; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5510 => 			--11
	if (mulfprdy = '1') then state := s5511;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5510; end if;
when s5511 => state := s5512; 	--12
	mulfpsclr <= '0';
when s5512 => state := s5513; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5513 => 			--14
	if (addfprdy = '1') then state := s5514;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5513; end if;
when s5514 => state := s5515; 	--15
	addfpsclr <= '0';
when s5515 => state := s5516; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5516 => 			--17
	if (addfprdy = '1') then state := s5517;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5516; end if;
when s5517 => state := s5518; 	--18
	addfpsclr <= '0';
when s5518 => state := s5519; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5519 => 			--20
	if (addfprdy = '1') then state := s5520;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5519; end if;
when s5520 => state := s5521; 	--21
	addfpsclr <= '0';
when s5521 => state := s5522; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (306, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5522 => state := s5523; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (550, 12)); -- offset LSB 502
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s5523 => state := s5524;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (551, 12)); -- offset MSB 503
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5524 => state := s5525; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5525 => 			--4
	if (fixed2floatrdy = '1') then state := s5526;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5525; end if;
when s5526 => state := s5527; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5527 => 			--6
	if (mulfprdy = '1') then state := s5528;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5527; end if;
when s5528 => state := s5529; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5529 => 			--8
	if (mulfprdy = '1') then state := s5530;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5529; end if;
when s5530 => state := s5531; 	--9
	mulfpsclr <= '0';
when s5531 => state := s5532; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5532 => 			--11
	if (mulfprdy = '1') then state := s5533;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5532; end if;
when s5533 => state := s5534; 	--12
	mulfpsclr <= '0';
when s5534 => state := s5535; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5535 => 			--14
	if (addfprdy = '1') then state := s5536;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5535; end if;
when s5536 => state := s5537; 	--15
	addfpsclr <= '0';
when s5537 => state := s5538; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5538 => 			--17
	if (addfprdy = '1') then state := s5539;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5538; end if;
when s5539 => state := s5540; 	--18
	addfpsclr <= '0';
when s5540 => state := s5541; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5541 => 			--20
	if (addfprdy = '1') then state := s5542;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5541; end if;
when s5542 => state := s5543; 	--21
	addfpsclr <= '0';
when s5543 => state := s5544; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (307, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5544 => state := s5545; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (552, 12)); -- offset LSB 504
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s5545 => state := s5546;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (553, 12)); -- offset MSB 505
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5546 => state := s5547; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5547 => 			--4
	if (fixed2floatrdy = '1') then state := s5548;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5547; end if;
when s5548 => state := s5549; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5549 => 			--6
	if (mulfprdy = '1') then state := s5550;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5549; end if;
when s5550 => state := s5551; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5551 => 			--8
	if (mulfprdy = '1') then state := s5552;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5551; end if;
when s5552 => state := s5553; 	--9
	mulfpsclr <= '0';
when s5553 => state := s5554; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5554 => 			--11
	if (mulfprdy = '1') then state := s5555;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5554; end if;
when s5555 => state := s5556; 	--12
	mulfpsclr <= '0';
when s5556 => state := s5557; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5557 => 			--14
	if (addfprdy = '1') then state := s5558;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5557; end if;
when s5558 => state := s5559; 	--15
	addfpsclr <= '0';
when s5559 => state := s5560; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5560 => 			--17
	if (addfprdy = '1') then state := s5561;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5560; end if;
when s5561 => state := s5562; 	--18
	addfpsclr <= '0';
when s5562 => state := s5563; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5563 => 			--20
	if (addfprdy = '1') then state := s5564;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5563; end if;
when s5564 => state := s5565; 	--21
	addfpsclr <= '0';
when s5565 => state := s5566; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (308, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5566 => state := s5567; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (554, 12)); -- offset LSB 506
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s5567 => state := s5568;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (555, 12)); -- offset MSB 507
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5568 => state := s5569; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5569 => 			--4
	if (fixed2floatrdy = '1') then state := s5570;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5569; end if;
when s5570 => state := s5571; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5571 => 			--6
	if (mulfprdy = '1') then state := s5572;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5571; end if;
when s5572 => state := s5573; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5573 => 			--8
	if (mulfprdy = '1') then state := s5574;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5573; end if;
when s5574 => state := s5575; 	--9
	mulfpsclr <= '0';
when s5575 => state := s5576; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5576 => 			--11
	if (mulfprdy = '1') then state := s5577;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5576; end if;
when s5577 => state := s5578; 	--12
	mulfpsclr <= '0';
when s5578 => state := s5579; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5579 => 			--14
	if (addfprdy = '1') then state := s5580;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5579; end if;
when s5580 => state := s5581; 	--15
	addfpsclr <= '0';
when s5581 => state := s5582; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5582 => 			--17
	if (addfprdy = '1') then state := s5583;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5582; end if;
when s5583 => state := s5584; 	--18
	addfpsclr <= '0';
when s5584 => state := s5585; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5585 => 			--20
	if (addfprdy = '1') then state := s5586;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5585; end if;
when s5586 => state := s5587; 	--21
	addfpsclr <= '0';
when s5587 => state := s5588; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (309, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5588 => state := s5589; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (556, 12)); -- offset LSB 508
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s5589 => state := s5590;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (557, 12)); -- offset MSB 509
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5590 => state := s5591; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5591 => 			--4
	if (fixed2floatrdy = '1') then state := s5592;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5591; end if;
when s5592 => state := s5593; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5593 => 			--6
	if (mulfprdy = '1') then state := s5594;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5593; end if;
when s5594 => state := s5595; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5595 => 			--8
	if (mulfprdy = '1') then state := s5596;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5595; end if;
when s5596 => state := s5597; 	--9
	mulfpsclr <= '0';
when s5597 => state := s5598; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5598 => 			--11
	if (mulfprdy = '1') then state := s5599;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5598; end if;
when s5599 => state := s5600; 	--12
	mulfpsclr <= '0';
when s5600 => state := s5601; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5601 => 			--14
	if (addfprdy = '1') then state := s5602;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5601; end if;
when s5602 => state := s5603; 	--15
	addfpsclr <= '0';
when s5603 => state := s5604; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5604 => 			--17
	if (addfprdy = '1') then state := s5605;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5604; end if;
when s5605 => state := s5606; 	--18
	addfpsclr <= '0';
when s5606 => state := s5607; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5607 => 			--20
	if (addfprdy = '1') then state := s5608;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5607; end if;
when s5608 => state := s5609; 	--21
	addfpsclr <= '0';
when s5609 => state := s5610; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (310, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5610 => state := s5611; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (558, 12)); -- offset LSB 510
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s5611 => state := s5612;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (559, 12)); -- offset MSB 511
	addra <= std_logic_vector (to_unsigned (7, 10)); -- OCCrowI 7
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5612 => state := s5613; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5613 => 			--4
	if (fixed2floatrdy = '1') then state := s5614;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5613; end if;
when s5614 => state := s5615; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5615 => 			--6
	if (mulfprdy = '1') then state := s5616;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5615; end if;
when s5616 => state := s5617; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5617 => 			--8
	if (mulfprdy = '1') then state := s5618;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5617; end if;
when s5618 => state := s5619; 	--9
	mulfpsclr <= '0';
when s5619 => state := s5620; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5620 => 			--11
	if (mulfprdy = '1') then state := s5621;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5620; end if;
when s5621 => state := s5622; 	--12
	mulfpsclr <= '0';
when s5622 => state := s5623; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5623 => 			--14
	if (addfprdy = '1') then state := s5624;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5623; end if;
when s5624 => state := s5625; 	--15
	addfpsclr <= '0';
when s5625 => state := s5626; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5626 => 			--17
	if (addfprdy = '1') then state := s5627;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5626; end if;
when s5627 => state := s5628; 	--18
	addfpsclr <= '0';
when s5628 => state := s5629; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5629 => 			--20
	if (addfprdy = '1') then state := s5630;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5629; end if;
when s5630 => state := s5631; 	--21
	addfpsclr <= '0';
when s5631 => state := s5632; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (311, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5632 => state := s5633; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (560, 12)); -- offset LSB 512
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s5633 => state := s5634;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (561, 12)); -- offset MSB 513
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5634 => state := s5635; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5635 => 			--4
	if (fixed2floatrdy = '1') then state := s5636;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5635; end if;
when s5636 => state := s5637; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5637 => 			--6
	if (mulfprdy = '1') then state := s5638;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5637; end if;
when s5638 => state := s5639; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5639 => 			--8
	if (mulfprdy = '1') then state := s5640;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5639; end if;
when s5640 => state := s5641; 	--9
	mulfpsclr <= '0';
when s5641 => state := s5642; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5642 => 			--11
	if (mulfprdy = '1') then state := s5643;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5642; end if;
when s5643 => state := s5644; 	--12
	mulfpsclr <= '0';
when s5644 => state := s5645; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5645 => 			--14
	if (addfprdy = '1') then state := s5646;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5645; end if;
when s5646 => state := s5647; 	--15
	addfpsclr <= '0';
when s5647 => state := s5648; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5648 => 			--17
	if (addfprdy = '1') then state := s5649;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5648; end if;
when s5649 => state := s5650; 	--18
	addfpsclr <= '0';
when s5650 => state := s5651; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5651 => 			--20
	if (addfprdy = '1') then state := s5652;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5651; end if;
when s5652 => state := s5653; 	--21
	addfpsclr <= '0';
when s5653 => state := s5654; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (312, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5654 => state := s5655; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (562, 12)); -- offset LSB 514
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s5655 => state := s5656;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (563, 12)); -- offset MSB 515
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5656 => state := s5657; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5657 => 			--4
	if (fixed2floatrdy = '1') then state := s5658;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5657; end if;
when s5658 => state := s5659; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5659 => 			--6
	if (mulfprdy = '1') then state := s5660;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5659; end if;
when s5660 => state := s5661; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5661 => 			--8
	if (mulfprdy = '1') then state := s5662;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5661; end if;
when s5662 => state := s5663; 	--9
	mulfpsclr <= '0';
when s5663 => state := s5664; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5664 => 			--11
	if (mulfprdy = '1') then state := s5665;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5664; end if;
when s5665 => state := s5666; 	--12
	mulfpsclr <= '0';
when s5666 => state := s5667; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5667 => 			--14
	if (addfprdy = '1') then state := s5668;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5667; end if;
when s5668 => state := s5669; 	--15
	addfpsclr <= '0';
when s5669 => state := s5670; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5670 => 			--17
	if (addfprdy = '1') then state := s5671;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5670; end if;
when s5671 => state := s5672; 	--18
	addfpsclr <= '0';
when s5672 => state := s5673; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5673 => 			--20
	if (addfprdy = '1') then state := s5674;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5673; end if;
when s5674 => state := s5675; 	--21
	addfpsclr <= '0';
when s5675 => state := s5676; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (313, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5676 => state := s5677; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (564, 12)); -- offset LSB 516
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s5677 => state := s5678;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (565, 12)); -- offset MSB 517
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5678 => state := s5679; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5679 => 			--4
	if (fixed2floatrdy = '1') then state := s5680;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5679; end if;
when s5680 => state := s5681; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5681 => 			--6
	if (mulfprdy = '1') then state := s5682;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5681; end if;
when s5682 => state := s5683; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5683 => 			--8
	if (mulfprdy = '1') then state := s5684;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5683; end if;
when s5684 => state := s5685; 	--9
	mulfpsclr <= '0';
when s5685 => state := s5686; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5686 => 			--11
	if (mulfprdy = '1') then state := s5687;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5686; end if;
when s5687 => state := s5688; 	--12
	mulfpsclr <= '0';
when s5688 => state := s5689; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5689 => 			--14
	if (addfprdy = '1') then state := s5690;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5689; end if;
when s5690 => state := s5691; 	--15
	addfpsclr <= '0';
when s5691 => state := s5692; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5692 => 			--17
	if (addfprdy = '1') then state := s5693;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5692; end if;
when s5693 => state := s5694; 	--18
	addfpsclr <= '0';
when s5694 => state := s5695; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5695 => 			--20
	if (addfprdy = '1') then state := s5696;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5695; end if;
when s5696 => state := s5697; 	--21
	addfpsclr <= '0';
when s5697 => state := s5698; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (314, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5698 => state := s5699; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (566, 12)); -- offset LSB 518
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s5699 => state := s5700;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (567, 12)); -- offset MSB 519
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5700 => state := s5701; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5701 => 			--4
	if (fixed2floatrdy = '1') then state := s5702;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5701; end if;
when s5702 => state := s5703; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5703 => 			--6
	if (mulfprdy = '1') then state := s5704;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5703; end if;
when s5704 => state := s5705; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5705 => 			--8
	if (mulfprdy = '1') then state := s5706;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5705; end if;
when s5706 => state := s5707; 	--9
	mulfpsclr <= '0';
when s5707 => state := s5708; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5708 => 			--11
	if (mulfprdy = '1') then state := s5709;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5708; end if;
when s5709 => state := s5710; 	--12
	mulfpsclr <= '0';
when s5710 => state := s5711; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5711 => 			--14
	if (addfprdy = '1') then state := s5712;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5711; end if;
when s5712 => state := s5713; 	--15
	addfpsclr <= '0';
when s5713 => state := s5714; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5714 => 			--17
	if (addfprdy = '1') then state := s5715;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5714; end if;
when s5715 => state := s5716; 	--18
	addfpsclr <= '0';
when s5716 => state := s5717; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5717 => 			--20
	if (addfprdy = '1') then state := s5718;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5717; end if;
when s5718 => state := s5719; 	--21
	addfpsclr <= '0';
when s5719 => state := s5720; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (315, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5720 => state := s5721; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (568, 12)); -- offset LSB 520
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s5721 => state := s5722;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (569, 12)); -- offset MSB 521
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5722 => state := s5723; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5723 => 			--4
	if (fixed2floatrdy = '1') then state := s5724;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5723; end if;
when s5724 => state := s5725; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5725 => 			--6
	if (mulfprdy = '1') then state := s5726;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5725; end if;
when s5726 => state := s5727; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5727 => 			--8
	if (mulfprdy = '1') then state := s5728;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5727; end if;
when s5728 => state := s5729; 	--9
	mulfpsclr <= '0';
when s5729 => state := s5730; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5730 => 			--11
	if (mulfprdy = '1') then state := s5731;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5730; end if;
when s5731 => state := s5732; 	--12
	mulfpsclr <= '0';
when s5732 => state := s5733; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5733 => 			--14
	if (addfprdy = '1') then state := s5734;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5733; end if;
when s5734 => state := s5735; 	--15
	addfpsclr <= '0';
when s5735 => state := s5736; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5736 => 			--17
	if (addfprdy = '1') then state := s5737;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5736; end if;
when s5737 => state := s5738; 	--18
	addfpsclr <= '0';
when s5738 => state := s5739; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5739 => 			--20
	if (addfprdy = '1') then state := s5740;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5739; end if;
when s5740 => state := s5741; 	--21
	addfpsclr <= '0';
when s5741 => state := s5742; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (316, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5742 => state := s5743; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (570, 12)); -- offset LSB 522
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s5743 => state := s5744;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (571, 12)); -- offset MSB 523
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5744 => state := s5745; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5745 => 			--4
	if (fixed2floatrdy = '1') then state := s5746;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5745; end if;
when s5746 => state := s5747; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5747 => 			--6
	if (mulfprdy = '1') then state := s5748;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5747; end if;
when s5748 => state := s5749; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5749 => 			--8
	if (mulfprdy = '1') then state := s5750;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5749; end if;
when s5750 => state := s5751; 	--9
	mulfpsclr <= '0';
when s5751 => state := s5752; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5752 => 			--11
	if (mulfprdy = '1') then state := s5753;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5752; end if;
when s5753 => state := s5754; 	--12
	mulfpsclr <= '0';
when s5754 => state := s5755; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5755 => 			--14
	if (addfprdy = '1') then state := s5756;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5755; end if;
when s5756 => state := s5757; 	--15
	addfpsclr <= '0';
when s5757 => state := s5758; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5758 => 			--17
	if (addfprdy = '1') then state := s5759;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5758; end if;
when s5759 => state := s5760; 	--18
	addfpsclr <= '0';
when s5760 => state := s5761; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5761 => 			--20
	if (addfprdy = '1') then state := s5762;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5761; end if;
when s5762 => state := s5763; 	--21
	addfpsclr <= '0';
when s5763 => state := s5764; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (317, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5764 => state := s5765; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (572, 12)); -- offset LSB 524
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s5765 => state := s5766;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (573, 12)); -- offset MSB 525
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5766 => state := s5767; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5767 => 			--4
	if (fixed2floatrdy = '1') then state := s5768;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5767; end if;
when s5768 => state := s5769; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5769 => 			--6
	if (mulfprdy = '1') then state := s5770;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5769; end if;
when s5770 => state := s5771; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5771 => 			--8
	if (mulfprdy = '1') then state := s5772;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5771; end if;
when s5772 => state := s5773; 	--9
	mulfpsclr <= '0';
when s5773 => state := s5774; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5774 => 			--11
	if (mulfprdy = '1') then state := s5775;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5774; end if;
when s5775 => state := s5776; 	--12
	mulfpsclr <= '0';
when s5776 => state := s5777; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5777 => 			--14
	if (addfprdy = '1') then state := s5778;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5777; end if;
when s5778 => state := s5779; 	--15
	addfpsclr <= '0';
when s5779 => state := s5780; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5780 => 			--17
	if (addfprdy = '1') then state := s5781;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5780; end if;
when s5781 => state := s5782; 	--18
	addfpsclr <= '0';
when s5782 => state := s5783; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5783 => 			--20
	if (addfprdy = '1') then state := s5784;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5783; end if;
when s5784 => state := s5785; 	--21
	addfpsclr <= '0';
when s5785 => state := s5786; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (318, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5786 => state := s5787; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (574, 12)); -- offset LSB 526
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s5787 => state := s5788;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (575, 12)); -- offset MSB 527
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5788 => state := s5789; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5789 => 			--4
	if (fixed2floatrdy = '1') then state := s5790;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5789; end if;
when s5790 => state := s5791; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5791 => 			--6
	if (mulfprdy = '1') then state := s5792;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5791; end if;
when s5792 => state := s5793; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5793 => 			--8
	if (mulfprdy = '1') then state := s5794;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5793; end if;
when s5794 => state := s5795; 	--9
	mulfpsclr <= '0';
when s5795 => state := s5796; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5796 => 			--11
	if (mulfprdy = '1') then state := s5797;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5796; end if;
when s5797 => state := s5798; 	--12
	mulfpsclr <= '0';
when s5798 => state := s5799; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5799 => 			--14
	if (addfprdy = '1') then state := s5800;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5799; end if;
when s5800 => state := s5801; 	--15
	addfpsclr <= '0';
when s5801 => state := s5802; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5802 => 			--17
	if (addfprdy = '1') then state := s5803;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5802; end if;
when s5803 => state := s5804; 	--18
	addfpsclr <= '0';
when s5804 => state := s5805; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5805 => 			--20
	if (addfprdy = '1') then state := s5806;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5805; end if;
when s5806 => state := s5807; 	--21
	addfpsclr <= '0';
when s5807 => state := s5808; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (319, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5808 => state := s5809; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (576, 12)); -- offset LSB 528
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s5809 => state := s5810;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (577, 12)); -- offset MSB 529
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5810 => state := s5811; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5811 => 			--4
	if (fixed2floatrdy = '1') then state := s5812;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5811; end if;
when s5812 => state := s5813; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5813 => 			--6
	if (mulfprdy = '1') then state := s5814;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5813; end if;
when s5814 => state := s5815; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5815 => 			--8
	if (mulfprdy = '1') then state := s5816;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5815; end if;
when s5816 => state := s5817; 	--9
	mulfpsclr <= '0';
when s5817 => state := s5818; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5818 => 			--11
	if (mulfprdy = '1') then state := s5819;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5818; end if;
when s5819 => state := s5820; 	--12
	mulfpsclr <= '0';
when s5820 => state := s5821; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5821 => 			--14
	if (addfprdy = '1') then state := s5822;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5821; end if;
when s5822 => state := s5823; 	--15
	addfpsclr <= '0';
when s5823 => state := s5824; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5824 => 			--17
	if (addfprdy = '1') then state := s5825;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5824; end if;
when s5825 => state := s5826; 	--18
	addfpsclr <= '0';
when s5826 => state := s5827; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5827 => 			--20
	if (addfprdy = '1') then state := s5828;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5827; end if;
when s5828 => state := s5829; 	--21
	addfpsclr <= '0';
when s5829 => state := s5830; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (320, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5830 => state := s5831; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (578, 12)); -- offset LSB 530
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s5831 => state := s5832;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (579, 12)); -- offset MSB 531
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5832 => state := s5833; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5833 => 			--4
	if (fixed2floatrdy = '1') then state := s5834;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5833; end if;
when s5834 => state := s5835; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5835 => 			--6
	if (mulfprdy = '1') then state := s5836;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5835; end if;
when s5836 => state := s5837; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5837 => 			--8
	if (mulfprdy = '1') then state := s5838;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5837; end if;
when s5838 => state := s5839; 	--9
	mulfpsclr <= '0';
when s5839 => state := s5840; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5840 => 			--11
	if (mulfprdy = '1') then state := s5841;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5840; end if;
when s5841 => state := s5842; 	--12
	mulfpsclr <= '0';
when s5842 => state := s5843; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5843 => 			--14
	if (addfprdy = '1') then state := s5844;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5843; end if;
when s5844 => state := s5845; 	--15
	addfpsclr <= '0';
when s5845 => state := s5846; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5846 => 			--17
	if (addfprdy = '1') then state := s5847;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5846; end if;
when s5847 => state := s5848; 	--18
	addfpsclr <= '0';
when s5848 => state := s5849; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5849 => 			--20
	if (addfprdy = '1') then state := s5850;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5849; end if;
when s5850 => state := s5851; 	--21
	addfpsclr <= '0';
when s5851 => state := s5852; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (321, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5852 => state := s5853; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (580, 12)); -- offset LSB 532
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s5853 => state := s5854;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (581, 12)); -- offset MSB 533
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5854 => state := s5855; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5855 => 			--4
	if (fixed2floatrdy = '1') then state := s5856;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5855; end if;
when s5856 => state := s5857; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5857 => 			--6
	if (mulfprdy = '1') then state := s5858;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5857; end if;
when s5858 => state := s5859; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5859 => 			--8
	if (mulfprdy = '1') then state := s5860;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5859; end if;
when s5860 => state := s5861; 	--9
	mulfpsclr <= '0';
when s5861 => state := s5862; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5862 => 			--11
	if (mulfprdy = '1') then state := s5863;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5862; end if;
when s5863 => state := s5864; 	--12
	mulfpsclr <= '0';
when s5864 => state := s5865; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5865 => 			--14
	if (addfprdy = '1') then state := s5866;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5865; end if;
when s5866 => state := s5867; 	--15
	addfpsclr <= '0';
when s5867 => state := s5868; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5868 => 			--17
	if (addfprdy = '1') then state := s5869;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5868; end if;
when s5869 => state := s5870; 	--18
	addfpsclr <= '0';
when s5870 => state := s5871; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5871 => 			--20
	if (addfprdy = '1') then state := s5872;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5871; end if;
when s5872 => state := s5873; 	--21
	addfpsclr <= '0';
when s5873 => state := s5874; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (322, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5874 => state := s5875; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (582, 12)); -- offset LSB 534
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s5875 => state := s5876;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (583, 12)); -- offset MSB 535
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5876 => state := s5877; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5877 => 			--4
	if (fixed2floatrdy = '1') then state := s5878;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5877; end if;
when s5878 => state := s5879; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5879 => 			--6
	if (mulfprdy = '1') then state := s5880;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5879; end if;
when s5880 => state := s5881; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5881 => 			--8
	if (mulfprdy = '1') then state := s5882;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5881; end if;
when s5882 => state := s5883; 	--9
	mulfpsclr <= '0';
when s5883 => state := s5884; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5884 => 			--11
	if (mulfprdy = '1') then state := s5885;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5884; end if;
when s5885 => state := s5886; 	--12
	mulfpsclr <= '0';
when s5886 => state := s5887; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5887 => 			--14
	if (addfprdy = '1') then state := s5888;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5887; end if;
when s5888 => state := s5889; 	--15
	addfpsclr <= '0';
when s5889 => state := s5890; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5890 => 			--17
	if (addfprdy = '1') then state := s5891;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5890; end if;
when s5891 => state := s5892; 	--18
	addfpsclr <= '0';
when s5892 => state := s5893; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5893 => 			--20
	if (addfprdy = '1') then state := s5894;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5893; end if;
when s5894 => state := s5895; 	--21
	addfpsclr <= '0';
when s5895 => state := s5896; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (323, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5896 => state := s5897; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (584, 12)); -- offset LSB 536
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s5897 => state := s5898;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (585, 12)); -- offset MSB 537
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5898 => state := s5899; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5899 => 			--4
	if (fixed2floatrdy = '1') then state := s5900;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5899; end if;
when s5900 => state := s5901; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5901 => 			--6
	if (mulfprdy = '1') then state := s5902;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5901; end if;
when s5902 => state := s5903; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5903 => 			--8
	if (mulfprdy = '1') then state := s5904;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5903; end if;
when s5904 => state := s5905; 	--9
	mulfpsclr <= '0';
when s5905 => state := s5906; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5906 => 			--11
	if (mulfprdy = '1') then state := s5907;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5906; end if;
when s5907 => state := s5908; 	--12
	mulfpsclr <= '0';
when s5908 => state := s5909; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5909 => 			--14
	if (addfprdy = '1') then state := s5910;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5909; end if;
when s5910 => state := s5911; 	--15
	addfpsclr <= '0';
when s5911 => state := s5912; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5912 => 			--17
	if (addfprdy = '1') then state := s5913;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5912; end if;
when s5913 => state := s5914; 	--18
	addfpsclr <= '0';
when s5914 => state := s5915; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5915 => 			--20
	if (addfprdy = '1') then state := s5916;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5915; end if;
when s5916 => state := s5917; 	--21
	addfpsclr <= '0';
when s5917 => state := s5918; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (324, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5918 => state := s5919; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (586, 12)); -- offset LSB 538
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s5919 => state := s5920;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (587, 12)); -- offset MSB 539
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5920 => state := s5921; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5921 => 			--4
	if (fixed2floatrdy = '1') then state := s5922;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5921; end if;
when s5922 => state := s5923; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5923 => 			--6
	if (mulfprdy = '1') then state := s5924;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5923; end if;
when s5924 => state := s5925; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5925 => 			--8
	if (mulfprdy = '1') then state := s5926;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5925; end if;
when s5926 => state := s5927; 	--9
	mulfpsclr <= '0';
when s5927 => state := s5928; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5928 => 			--11
	if (mulfprdy = '1') then state := s5929;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5928; end if;
when s5929 => state := s5930; 	--12
	mulfpsclr <= '0';
when s5930 => state := s5931; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5931 => 			--14
	if (addfprdy = '1') then state := s5932;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5931; end if;
when s5932 => state := s5933; 	--15
	addfpsclr <= '0';
when s5933 => state := s5934; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5934 => 			--17
	if (addfprdy = '1') then state := s5935;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5934; end if;
when s5935 => state := s5936; 	--18
	addfpsclr <= '0';
when s5936 => state := s5937; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5937 => 			--20
	if (addfprdy = '1') then state := s5938;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5937; end if;
when s5938 => state := s5939; 	--21
	addfpsclr <= '0';
when s5939 => state := s5940; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (325, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5940 => state := s5941; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (588, 12)); -- offset LSB 540
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s5941 => state := s5942;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (589, 12)); -- offset MSB 541
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5942 => state := s5943; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5943 => 			--4
	if (fixed2floatrdy = '1') then state := s5944;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5943; end if;
when s5944 => state := s5945; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5945 => 			--6
	if (mulfprdy = '1') then state := s5946;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5945; end if;
when s5946 => state := s5947; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5947 => 			--8
	if (mulfprdy = '1') then state := s5948;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5947; end if;
when s5948 => state := s5949; 	--9
	mulfpsclr <= '0';
when s5949 => state := s5950; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5950 => 			--11
	if (mulfprdy = '1') then state := s5951;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5950; end if;
when s5951 => state := s5952; 	--12
	mulfpsclr <= '0';
when s5952 => state := s5953; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5953 => 			--14
	if (addfprdy = '1') then state := s5954;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5953; end if;
when s5954 => state := s5955; 	--15
	addfpsclr <= '0';
when s5955 => state := s5956; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5956 => 			--17
	if (addfprdy = '1') then state := s5957;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5956; end if;
when s5957 => state := s5958; 	--18
	addfpsclr <= '0';
when s5958 => state := s5959; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5959 => 			--20
	if (addfprdy = '1') then state := s5960;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5959; end if;
when s5960 => state := s5961; 	--21
	addfpsclr <= '0';
when s5961 => state := s5962; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (326, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5962 => state := s5963; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (590, 12)); -- offset LSB 542
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s5963 => state := s5964;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (591, 12)); -- offset MSB 543
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5964 => state := s5965; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5965 => 			--4
	if (fixed2floatrdy = '1') then state := s5966;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5965; end if;
when s5966 => state := s5967; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5967 => 			--6
	if (mulfprdy = '1') then state := s5968;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5967; end if;
when s5968 => state := s5969; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5969 => 			--8
	if (mulfprdy = '1') then state := s5970;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5969; end if;
when s5970 => state := s5971; 	--9
	mulfpsclr <= '0';
when s5971 => state := s5972; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5972 => 			--11
	if (mulfprdy = '1') then state := s5973;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5972; end if;
when s5973 => state := s5974; 	--12
	mulfpsclr <= '0';
when s5974 => state := s5975; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5975 => 			--14
	if (addfprdy = '1') then state := s5976;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5975; end if;
when s5976 => state := s5977; 	--15
	addfpsclr <= '0';
when s5977 => state := s5978; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s5978 => 			--17
	if (addfprdy = '1') then state := s5979;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5978; end if;
when s5979 => state := s5980; 	--18
	addfpsclr <= '0';
when s5980 => state := s5981; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s5981 => 			--20
	if (addfprdy = '1') then state := s5982;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5981; end if;
when s5982 => state := s5983; 	--21
	addfpsclr <= '0';
when s5983 => state := s5984; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (327, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s5984 => state := s5985; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (592, 12)); -- offset LSB 544
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s5985 => state := s5986;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (593, 12)); -- offset MSB 545
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s5986 => state := s5987; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s5987 => 			--4
	if (fixed2floatrdy = '1') then state := s5988;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s5987; end if;
when s5988 => state := s5989; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s5989 => 			--6
	if (mulfprdy = '1') then state := s5990;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5989; end if;
when s5990 => state := s5991; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s5991 => 			--8
	if (mulfprdy = '1') then state := s5992;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5991; end if;
when s5992 => state := s5993; 	--9
	mulfpsclr <= '0';
when s5993 => state := s5994; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s5994 => 			--11
	if (mulfprdy = '1') then state := s5995;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s5994; end if;
when s5995 => state := s5996; 	--12
	mulfpsclr <= '0';
when s5996 => state := s5997; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s5997 => 			--14
	if (addfprdy = '1') then state := s5998;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s5997; end if;
when s5998 => state := s5999; 	--15
	addfpsclr <= '0';
when s5999 => state := s6000; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6000 => 			--17
	if (addfprdy = '1') then state := s6001;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6000; end if;
when s6001 => state := s6002; 	--18
	addfpsclr <= '0';
when s6002 => state := s6003; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6003 => 			--20
	if (addfprdy = '1') then state := s6004;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6003; end if;
when s6004 => state := s6005; 	--21
	addfpsclr <= '0';
when s6005 => state := s6006; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (328, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6006 => state := s6007; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (594, 12)); -- offset LSB 546
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s6007 => state := s6008;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (595, 12)); -- offset MSB 547
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6008 => state := s6009; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6009 => 			--4
	if (fixed2floatrdy = '1') then state := s6010;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6009; end if;
when s6010 => state := s6011; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6011 => 			--6
	if (mulfprdy = '1') then state := s6012;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6011; end if;
when s6012 => state := s6013; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6013 => 			--8
	if (mulfprdy = '1') then state := s6014;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6013; end if;
when s6014 => state := s6015; 	--9
	mulfpsclr <= '0';
when s6015 => state := s6016; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6016 => 			--11
	if (mulfprdy = '1') then state := s6017;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6016; end if;
when s6017 => state := s6018; 	--12
	mulfpsclr <= '0';
when s6018 => state := s6019; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6019 => 			--14
	if (addfprdy = '1') then state := s6020;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6019; end if;
when s6020 => state := s6021; 	--15
	addfpsclr <= '0';
when s6021 => state := s6022; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6022 => 			--17
	if (addfprdy = '1') then state := s6023;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6022; end if;
when s6023 => state := s6024; 	--18
	addfpsclr <= '0';
when s6024 => state := s6025; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6025 => 			--20
	if (addfprdy = '1') then state := s6026;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6025; end if;
when s6026 => state := s6027; 	--21
	addfpsclr <= '0';
when s6027 => state := s6028; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (329, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6028 => state := s6029; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (596, 12)); -- offset LSB 548
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s6029 => state := s6030;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (597, 12)); -- offset MSB 549
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6030 => state := s6031; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6031 => 			--4
	if (fixed2floatrdy = '1') then state := s6032;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6031; end if;
when s6032 => state := s6033; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6033 => 			--6
	if (mulfprdy = '1') then state := s6034;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6033; end if;
when s6034 => state := s6035; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6035 => 			--8
	if (mulfprdy = '1') then state := s6036;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6035; end if;
when s6036 => state := s6037; 	--9
	mulfpsclr <= '0';
when s6037 => state := s6038; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6038 => 			--11
	if (mulfprdy = '1') then state := s6039;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6038; end if;
when s6039 => state := s6040; 	--12
	mulfpsclr <= '0';
when s6040 => state := s6041; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6041 => 			--14
	if (addfprdy = '1') then state := s6042;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6041; end if;
when s6042 => state := s6043; 	--15
	addfpsclr <= '0';
when s6043 => state := s6044; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6044 => 			--17
	if (addfprdy = '1') then state := s6045;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6044; end if;
when s6045 => state := s6046; 	--18
	addfpsclr <= '0';
when s6046 => state := s6047; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6047 => 			--20
	if (addfprdy = '1') then state := s6048;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6047; end if;
when s6048 => state := s6049; 	--21
	addfpsclr <= '0';
when s6049 => state := s6050; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (330, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6050 => state := s6051; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (598, 12)); -- offset LSB 550
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s6051 => state := s6052;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (599, 12)); -- offset MSB 551
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6052 => state := s6053; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6053 => 			--4
	if (fixed2floatrdy = '1') then state := s6054;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6053; end if;
when s6054 => state := s6055; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6055 => 			--6
	if (mulfprdy = '1') then state := s6056;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6055; end if;
when s6056 => state := s6057; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6057 => 			--8
	if (mulfprdy = '1') then state := s6058;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6057; end if;
when s6058 => state := s6059; 	--9
	mulfpsclr <= '0';
when s6059 => state := s6060; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6060 => 			--11
	if (mulfprdy = '1') then state := s6061;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6060; end if;
when s6061 => state := s6062; 	--12
	mulfpsclr <= '0';
when s6062 => state := s6063; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6063 => 			--14
	if (addfprdy = '1') then state := s6064;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6063; end if;
when s6064 => state := s6065; 	--15
	addfpsclr <= '0';
when s6065 => state := s6066; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6066 => 			--17
	if (addfprdy = '1') then state := s6067;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6066; end if;
when s6067 => state := s6068; 	--18
	addfpsclr <= '0';
when s6068 => state := s6069; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6069 => 			--20
	if (addfprdy = '1') then state := s6070;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6069; end if;
when s6070 => state := s6071; 	--21
	addfpsclr <= '0';
when s6071 => state := s6072; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (331, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6072 => state := s6073; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (600, 12)); -- offset LSB 552
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s6073 => state := s6074;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (601, 12)); -- offset MSB 553
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6074 => state := s6075; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6075 => 			--4
	if (fixed2floatrdy = '1') then state := s6076;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6075; end if;
when s6076 => state := s6077; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6077 => 			--6
	if (mulfprdy = '1') then state := s6078;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6077; end if;
when s6078 => state := s6079; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6079 => 			--8
	if (mulfprdy = '1') then state := s6080;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6079; end if;
when s6080 => state := s6081; 	--9
	mulfpsclr <= '0';
when s6081 => state := s6082; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6082 => 			--11
	if (mulfprdy = '1') then state := s6083;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6082; end if;
when s6083 => state := s6084; 	--12
	mulfpsclr <= '0';
when s6084 => state := s6085; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6085 => 			--14
	if (addfprdy = '1') then state := s6086;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6085; end if;
when s6086 => state := s6087; 	--15
	addfpsclr <= '0';
when s6087 => state := s6088; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6088 => 			--17
	if (addfprdy = '1') then state := s6089;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6088; end if;
when s6089 => state := s6090; 	--18
	addfpsclr <= '0';
when s6090 => state := s6091; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6091 => 			--20
	if (addfprdy = '1') then state := s6092;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6091; end if;
when s6092 => state := s6093; 	--21
	addfpsclr <= '0';
when s6093 => state := s6094; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (332, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6094 => state := s6095; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (602, 12)); -- offset LSB 554
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s6095 => state := s6096;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (603, 12)); -- offset MSB 555
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6096 => state := s6097; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6097 => 			--4
	if (fixed2floatrdy = '1') then state := s6098;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6097; end if;
when s6098 => state := s6099; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6099 => 			--6
	if (mulfprdy = '1') then state := s6100;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6099; end if;
when s6100 => state := s6101; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6101 => 			--8
	if (mulfprdy = '1') then state := s6102;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6101; end if;
when s6102 => state := s6103; 	--9
	mulfpsclr <= '0';
when s6103 => state := s6104; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6104 => 			--11
	if (mulfprdy = '1') then state := s6105;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6104; end if;
when s6105 => state := s6106; 	--12
	mulfpsclr <= '0';
when s6106 => state := s6107; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6107 => 			--14
	if (addfprdy = '1') then state := s6108;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6107; end if;
when s6108 => state := s6109; 	--15
	addfpsclr <= '0';
when s6109 => state := s6110; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6110 => 			--17
	if (addfprdy = '1') then state := s6111;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6110; end if;
when s6111 => state := s6112; 	--18
	addfpsclr <= '0';
when s6112 => state := s6113; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6113 => 			--20
	if (addfprdy = '1') then state := s6114;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6113; end if;
when s6114 => state := s6115; 	--21
	addfpsclr <= '0';
when s6115 => state := s6116; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (333, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6116 => state := s6117; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (604, 12)); -- offset LSB 556
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s6117 => state := s6118;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (605, 12)); -- offset MSB 557
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6118 => state := s6119; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6119 => 			--4
	if (fixed2floatrdy = '1') then state := s6120;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6119; end if;
when s6120 => state := s6121; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6121 => 			--6
	if (mulfprdy = '1') then state := s6122;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6121; end if;
when s6122 => state := s6123; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6123 => 			--8
	if (mulfprdy = '1') then state := s6124;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6123; end if;
when s6124 => state := s6125; 	--9
	mulfpsclr <= '0';
when s6125 => state := s6126; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6126 => 			--11
	if (mulfprdy = '1') then state := s6127;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6126; end if;
when s6127 => state := s6128; 	--12
	mulfpsclr <= '0';
when s6128 => state := s6129; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6129 => 			--14
	if (addfprdy = '1') then state := s6130;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6129; end if;
when s6130 => state := s6131; 	--15
	addfpsclr <= '0';
when s6131 => state := s6132; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6132 => 			--17
	if (addfprdy = '1') then state := s6133;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6132; end if;
when s6133 => state := s6134; 	--18
	addfpsclr <= '0';
when s6134 => state := s6135; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6135 => 			--20
	if (addfprdy = '1') then state := s6136;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6135; end if;
when s6136 => state := s6137; 	--21
	addfpsclr <= '0';
when s6137 => state := s6138; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (334, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6138 => state := s6139; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (606, 12)); -- offset LSB 558
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s6139 => state := s6140;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (607, 12)); -- offset MSB 559
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6140 => state := s6141; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6141 => 			--4
	if (fixed2floatrdy = '1') then state := s6142;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6141; end if;
when s6142 => state := s6143; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6143 => 			--6
	if (mulfprdy = '1') then state := s6144;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6143; end if;
when s6144 => state := s6145; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6145 => 			--8
	if (mulfprdy = '1') then state := s6146;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6145; end if;
when s6146 => state := s6147; 	--9
	mulfpsclr <= '0';
when s6147 => state := s6148; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6148 => 			--11
	if (mulfprdy = '1') then state := s6149;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6148; end if;
when s6149 => state := s6150; 	--12
	mulfpsclr <= '0';
when s6150 => state := s6151; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6151 => 			--14
	if (addfprdy = '1') then state := s6152;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6151; end if;
when s6152 => state := s6153; 	--15
	addfpsclr <= '0';
when s6153 => state := s6154; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6154 => 			--17
	if (addfprdy = '1') then state := s6155;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6154; end if;
when s6155 => state := s6156; 	--18
	addfpsclr <= '0';
when s6156 => state := s6157; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6157 => 			--20
	if (addfprdy = '1') then state := s6158;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6157; end if;
when s6158 => state := s6159; 	--21
	addfpsclr <= '0';
when s6159 => state := s6160; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (335, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6160 => state := s6161; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (608, 12)); -- offset LSB 560
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s6161 => state := s6162;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (609, 12)); -- offset MSB 561
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6162 => state := s6163; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6163 => 			--4
	if (fixed2floatrdy = '1') then state := s6164;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6163; end if;
when s6164 => state := s6165; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6165 => 			--6
	if (mulfprdy = '1') then state := s6166;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6165; end if;
when s6166 => state := s6167; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6167 => 			--8
	if (mulfprdy = '1') then state := s6168;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6167; end if;
when s6168 => state := s6169; 	--9
	mulfpsclr <= '0';
when s6169 => state := s6170; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6170 => 			--11
	if (mulfprdy = '1') then state := s6171;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6170; end if;
when s6171 => state := s6172; 	--12
	mulfpsclr <= '0';
when s6172 => state := s6173; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6173 => 			--14
	if (addfprdy = '1') then state := s6174;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6173; end if;
when s6174 => state := s6175; 	--15
	addfpsclr <= '0';
when s6175 => state := s6176; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6176 => 			--17
	if (addfprdy = '1') then state := s6177;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6176; end if;
when s6177 => state := s6178; 	--18
	addfpsclr <= '0';
when s6178 => state := s6179; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6179 => 			--20
	if (addfprdy = '1') then state := s6180;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6179; end if;
when s6180 => state := s6181; 	--21
	addfpsclr <= '0';
when s6181 => state := s6182; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (336, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6182 => state := s6183; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (610, 12)); -- offset LSB 562
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s6183 => state := s6184;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (611, 12)); -- offset MSB 563
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6184 => state := s6185; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6185 => 			--4
	if (fixed2floatrdy = '1') then state := s6186;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6185; end if;
when s6186 => state := s6187; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6187 => 			--6
	if (mulfprdy = '1') then state := s6188;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6187; end if;
when s6188 => state := s6189; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6189 => 			--8
	if (mulfprdy = '1') then state := s6190;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6189; end if;
when s6190 => state := s6191; 	--9
	mulfpsclr <= '0';
when s6191 => state := s6192; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6192 => 			--11
	if (mulfprdy = '1') then state := s6193;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6192; end if;
when s6193 => state := s6194; 	--12
	mulfpsclr <= '0';
when s6194 => state := s6195; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6195 => 			--14
	if (addfprdy = '1') then state := s6196;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6195; end if;
when s6196 => state := s6197; 	--15
	addfpsclr <= '0';
when s6197 => state := s6198; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6198 => 			--17
	if (addfprdy = '1') then state := s6199;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6198; end if;
when s6199 => state := s6200; 	--18
	addfpsclr <= '0';
when s6200 => state := s6201; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6201 => 			--20
	if (addfprdy = '1') then state := s6202;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6201; end if;
when s6202 => state := s6203; 	--21
	addfpsclr <= '0';
when s6203 => state := s6204; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (337, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6204 => state := s6205; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (612, 12)); -- offset LSB 564
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s6205 => state := s6206;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (613, 12)); -- offset MSB 565
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6206 => state := s6207; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6207 => 			--4
	if (fixed2floatrdy = '1') then state := s6208;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6207; end if;
when s6208 => state := s6209; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6209 => 			--6
	if (mulfprdy = '1') then state := s6210;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6209; end if;
when s6210 => state := s6211; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6211 => 			--8
	if (mulfprdy = '1') then state := s6212;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6211; end if;
when s6212 => state := s6213; 	--9
	mulfpsclr <= '0';
when s6213 => state := s6214; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6214 => 			--11
	if (mulfprdy = '1') then state := s6215;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6214; end if;
when s6215 => state := s6216; 	--12
	mulfpsclr <= '0';
when s6216 => state := s6217; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6217 => 			--14
	if (addfprdy = '1') then state := s6218;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6217; end if;
when s6218 => state := s6219; 	--15
	addfpsclr <= '0';
when s6219 => state := s6220; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6220 => 			--17
	if (addfprdy = '1') then state := s6221;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6220; end if;
when s6221 => state := s6222; 	--18
	addfpsclr <= '0';
when s6222 => state := s6223; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6223 => 			--20
	if (addfprdy = '1') then state := s6224;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6223; end if;
when s6224 => state := s6225; 	--21
	addfpsclr <= '0';
when s6225 => state := s6226; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (338, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6226 => state := s6227; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (614, 12)); -- offset LSB 566
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s6227 => state := s6228;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (615, 12)); -- offset MSB 567
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6228 => state := s6229; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6229 => 			--4
	if (fixed2floatrdy = '1') then state := s6230;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6229; end if;
when s6230 => state := s6231; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6231 => 			--6
	if (mulfprdy = '1') then state := s6232;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6231; end if;
when s6232 => state := s6233; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6233 => 			--8
	if (mulfprdy = '1') then state := s6234;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6233; end if;
when s6234 => state := s6235; 	--9
	mulfpsclr <= '0';
when s6235 => state := s6236; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6236 => 			--11
	if (mulfprdy = '1') then state := s6237;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6236; end if;
when s6237 => state := s6238; 	--12
	mulfpsclr <= '0';
when s6238 => state := s6239; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6239 => 			--14
	if (addfprdy = '1') then state := s6240;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6239; end if;
when s6240 => state := s6241; 	--15
	addfpsclr <= '0';
when s6241 => state := s6242; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6242 => 			--17
	if (addfprdy = '1') then state := s6243;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6242; end if;
when s6243 => state := s6244; 	--18
	addfpsclr <= '0';
when s6244 => state := s6245; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6245 => 			--20
	if (addfprdy = '1') then state := s6246;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6245; end if;
when s6246 => state := s6247; 	--21
	addfpsclr <= '0';
when s6247 => state := s6248; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (339, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6248 => state := s6249; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (616, 12)); -- offset LSB 568
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s6249 => state := s6250;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (617, 12)); -- offset MSB 569
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6250 => state := s6251; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6251 => 			--4
	if (fixed2floatrdy = '1') then state := s6252;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6251; end if;
when s6252 => state := s6253; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6253 => 			--6
	if (mulfprdy = '1') then state := s6254;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6253; end if;
when s6254 => state := s6255; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6255 => 			--8
	if (mulfprdy = '1') then state := s6256;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6255; end if;
when s6256 => state := s6257; 	--9
	mulfpsclr <= '0';
when s6257 => state := s6258; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6258 => 			--11
	if (mulfprdy = '1') then state := s6259;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6258; end if;
when s6259 => state := s6260; 	--12
	mulfpsclr <= '0';
when s6260 => state := s6261; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6261 => 			--14
	if (addfprdy = '1') then state := s6262;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6261; end if;
when s6262 => state := s6263; 	--15
	addfpsclr <= '0';
when s6263 => state := s6264; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6264 => 			--17
	if (addfprdy = '1') then state := s6265;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6264; end if;
when s6265 => state := s6266; 	--18
	addfpsclr <= '0';
when s6266 => state := s6267; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6267 => 			--20
	if (addfprdy = '1') then state := s6268;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6267; end if;
when s6268 => state := s6269; 	--21
	addfpsclr <= '0';
when s6269 => state := s6270; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (340, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6270 => state := s6271; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (618, 12)); -- offset LSB 570
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s6271 => state := s6272;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (619, 12)); -- offset MSB 571
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6272 => state := s6273; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6273 => 			--4
	if (fixed2floatrdy = '1') then state := s6274;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6273; end if;
when s6274 => state := s6275; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6275 => 			--6
	if (mulfprdy = '1') then state := s6276;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6275; end if;
when s6276 => state := s6277; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6277 => 			--8
	if (mulfprdy = '1') then state := s6278;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6277; end if;
when s6278 => state := s6279; 	--9
	mulfpsclr <= '0';
when s6279 => state := s6280; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6280 => 			--11
	if (mulfprdy = '1') then state := s6281;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6280; end if;
when s6281 => state := s6282; 	--12
	mulfpsclr <= '0';
when s6282 => state := s6283; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6283 => 			--14
	if (addfprdy = '1') then state := s6284;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6283; end if;
when s6284 => state := s6285; 	--15
	addfpsclr <= '0';
when s6285 => state := s6286; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6286 => 			--17
	if (addfprdy = '1') then state := s6287;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6286; end if;
when s6287 => state := s6288; 	--18
	addfpsclr <= '0';
when s6288 => state := s6289; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6289 => 			--20
	if (addfprdy = '1') then state := s6290;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6289; end if;
when s6290 => state := s6291; 	--21
	addfpsclr <= '0';
when s6291 => state := s6292; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (341, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6292 => state := s6293; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (620, 12)); -- offset LSB 572
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s6293 => state := s6294;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (621, 12)); -- offset MSB 573
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6294 => state := s6295; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6295 => 			--4
	if (fixed2floatrdy = '1') then state := s6296;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6295; end if;
when s6296 => state := s6297; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6297 => 			--6
	if (mulfprdy = '1') then state := s6298;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6297; end if;
when s6298 => state := s6299; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6299 => 			--8
	if (mulfprdy = '1') then state := s6300;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6299; end if;
when s6300 => state := s6301; 	--9
	mulfpsclr <= '0';
when s6301 => state := s6302; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6302 => 			--11
	if (mulfprdy = '1') then state := s6303;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6302; end if;
when s6303 => state := s6304; 	--12
	mulfpsclr <= '0';
when s6304 => state := s6305; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6305 => 			--14
	if (addfprdy = '1') then state := s6306;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6305; end if;
when s6306 => state := s6307; 	--15
	addfpsclr <= '0';
when s6307 => state := s6308; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6308 => 			--17
	if (addfprdy = '1') then state := s6309;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6308; end if;
when s6309 => state := s6310; 	--18
	addfpsclr <= '0';
when s6310 => state := s6311; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6311 => 			--20
	if (addfprdy = '1') then state := s6312;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6311; end if;
when s6312 => state := s6313; 	--21
	addfpsclr <= '0';
when s6313 => state := s6314; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (342, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6314 => state := s6315; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (622, 12)); -- offset LSB 574
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s6315 => state := s6316;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (623, 12)); -- offset MSB 575
	addra <= std_logic_vector (to_unsigned (8, 10)); -- OCCrowI 8
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6316 => state := s6317; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6317 => 			--4
	if (fixed2floatrdy = '1') then state := s6318;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6317; end if;
when s6318 => state := s6319; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6319 => 			--6
	if (mulfprdy = '1') then state := s6320;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6319; end if;
when s6320 => state := s6321; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6321 => 			--8
	if (mulfprdy = '1') then state := s6322;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6321; end if;
when s6322 => state := s6323; 	--9
	mulfpsclr <= '0';
when s6323 => state := s6324; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6324 => 			--11
	if (mulfprdy = '1') then state := s6325;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6324; end if;
when s6325 => state := s6326; 	--12
	mulfpsclr <= '0';
when s6326 => state := s6327; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6327 => 			--14
	if (addfprdy = '1') then state := s6328;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6327; end if;
when s6328 => state := s6329; 	--15
	addfpsclr <= '0';
when s6329 => state := s6330; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6330 => 			--17
	if (addfprdy = '1') then state := s6331;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6330; end if;
when s6331 => state := s6332; 	--18
	addfpsclr <= '0';
when s6332 => state := s6333; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6333 => 			--20
	if (addfprdy = '1') then state := s6334;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6333; end if;
when s6334 => state := s6335; 	--21
	addfpsclr <= '0';
when s6335 => state := s6336; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (343, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6336 => state := s6337; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (624, 12)); -- offset LSB 576
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s6337 => state := s6338;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (625, 12)); -- offset MSB 577
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6338 => state := s6339; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6339 => 			--4
	if (fixed2floatrdy = '1') then state := s6340;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6339; end if;
when s6340 => state := s6341; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6341 => 			--6
	if (mulfprdy = '1') then state := s6342;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6341; end if;
when s6342 => state := s6343; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6343 => 			--8
	if (mulfprdy = '1') then state := s6344;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6343; end if;
when s6344 => state := s6345; 	--9
	mulfpsclr <= '0';
when s6345 => state := s6346; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6346 => 			--11
	if (mulfprdy = '1') then state := s6347;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6346; end if;
when s6347 => state := s6348; 	--12
	mulfpsclr <= '0';
when s6348 => state := s6349; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6349 => 			--14
	if (addfprdy = '1') then state := s6350;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6349; end if;
when s6350 => state := s6351; 	--15
	addfpsclr <= '0';
when s6351 => state := s6352; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6352 => 			--17
	if (addfprdy = '1') then state := s6353;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6352; end if;
when s6353 => state := s6354; 	--18
	addfpsclr <= '0';
when s6354 => state := s6355; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6355 => 			--20
	if (addfprdy = '1') then state := s6356;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6355; end if;
when s6356 => state := s6357; 	--21
	addfpsclr <= '0';
when s6357 => state := s6358; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (344, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6358 => state := s6359; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (626, 12)); -- offset LSB 578
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s6359 => state := s6360;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (627, 12)); -- offset MSB 579
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6360 => state := s6361; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6361 => 			--4
	if (fixed2floatrdy = '1') then state := s6362;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6361; end if;
when s6362 => state := s6363; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6363 => 			--6
	if (mulfprdy = '1') then state := s6364;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6363; end if;
when s6364 => state := s6365; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6365 => 			--8
	if (mulfprdy = '1') then state := s6366;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6365; end if;
when s6366 => state := s6367; 	--9
	mulfpsclr <= '0';
when s6367 => state := s6368; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6368 => 			--11
	if (mulfprdy = '1') then state := s6369;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6368; end if;
when s6369 => state := s6370; 	--12
	mulfpsclr <= '0';
when s6370 => state := s6371; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6371 => 			--14
	if (addfprdy = '1') then state := s6372;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6371; end if;
when s6372 => state := s6373; 	--15
	addfpsclr <= '0';
when s6373 => state := s6374; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6374 => 			--17
	if (addfprdy = '1') then state := s6375;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6374; end if;
when s6375 => state := s6376; 	--18
	addfpsclr <= '0';
when s6376 => state := s6377; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6377 => 			--20
	if (addfprdy = '1') then state := s6378;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6377; end if;
when s6378 => state := s6379; 	--21
	addfpsclr <= '0';
when s6379 => state := s6380; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (345, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6380 => state := s6381; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (628, 12)); -- offset LSB 580
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s6381 => state := s6382;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (629, 12)); -- offset MSB 581
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6382 => state := s6383; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6383 => 			--4
	if (fixed2floatrdy = '1') then state := s6384;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6383; end if;
when s6384 => state := s6385; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6385 => 			--6
	if (mulfprdy = '1') then state := s6386;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6385; end if;
when s6386 => state := s6387; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6387 => 			--8
	if (mulfprdy = '1') then state := s6388;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6387; end if;
when s6388 => state := s6389; 	--9
	mulfpsclr <= '0';
when s6389 => state := s6390; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6390 => 			--11
	if (mulfprdy = '1') then state := s6391;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6390; end if;
when s6391 => state := s6392; 	--12
	mulfpsclr <= '0';
when s6392 => state := s6393; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6393 => 			--14
	if (addfprdy = '1') then state := s6394;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6393; end if;
when s6394 => state := s6395; 	--15
	addfpsclr <= '0';
when s6395 => state := s6396; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6396 => 			--17
	if (addfprdy = '1') then state := s6397;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6396; end if;
when s6397 => state := s6398; 	--18
	addfpsclr <= '0';
when s6398 => state := s6399; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6399 => 			--20
	if (addfprdy = '1') then state := s6400;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6399; end if;
when s6400 => state := s6401; 	--21
	addfpsclr <= '0';
when s6401 => state := s6402; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (346, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6402 => state := s6403; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (630, 12)); -- offset LSB 582
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s6403 => state := s6404;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (631, 12)); -- offset MSB 583
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6404 => state := s6405; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6405 => 			--4
	if (fixed2floatrdy = '1') then state := s6406;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6405; end if;
when s6406 => state := s6407; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6407 => 			--6
	if (mulfprdy = '1') then state := s6408;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6407; end if;
when s6408 => state := s6409; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6409 => 			--8
	if (mulfprdy = '1') then state := s6410;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6409; end if;
when s6410 => state := s6411; 	--9
	mulfpsclr <= '0';
when s6411 => state := s6412; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6412 => 			--11
	if (mulfprdy = '1') then state := s6413;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6412; end if;
when s6413 => state := s6414; 	--12
	mulfpsclr <= '0';
when s6414 => state := s6415; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6415 => 			--14
	if (addfprdy = '1') then state := s6416;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6415; end if;
when s6416 => state := s6417; 	--15
	addfpsclr <= '0';
when s6417 => state := s6418; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6418 => 			--17
	if (addfprdy = '1') then state := s6419;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6418; end if;
when s6419 => state := s6420; 	--18
	addfpsclr <= '0';
when s6420 => state := s6421; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6421 => 			--20
	if (addfprdy = '1') then state := s6422;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6421; end if;
when s6422 => state := s6423; 	--21
	addfpsclr <= '0';
when s6423 => state := s6424; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (347, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6424 => state := s6425; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (632, 12)); -- offset LSB 584
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s6425 => state := s6426;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (633, 12)); -- offset MSB 585
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6426 => state := s6427; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6427 => 			--4
	if (fixed2floatrdy = '1') then state := s6428;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6427; end if;
when s6428 => state := s6429; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6429 => 			--6
	if (mulfprdy = '1') then state := s6430;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6429; end if;
when s6430 => state := s6431; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6431 => 			--8
	if (mulfprdy = '1') then state := s6432;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6431; end if;
when s6432 => state := s6433; 	--9
	mulfpsclr <= '0';
when s6433 => state := s6434; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6434 => 			--11
	if (mulfprdy = '1') then state := s6435;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6434; end if;
when s6435 => state := s6436; 	--12
	mulfpsclr <= '0';
when s6436 => state := s6437; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6437 => 			--14
	if (addfprdy = '1') then state := s6438;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6437; end if;
when s6438 => state := s6439; 	--15
	addfpsclr <= '0';
when s6439 => state := s6440; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6440 => 			--17
	if (addfprdy = '1') then state := s6441;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6440; end if;
when s6441 => state := s6442; 	--18
	addfpsclr <= '0';
when s6442 => state := s6443; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6443 => 			--20
	if (addfprdy = '1') then state := s6444;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6443; end if;
when s6444 => state := s6445; 	--21
	addfpsclr <= '0';
when s6445 => state := s6446; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (348, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6446 => state := s6447; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (634, 12)); -- offset LSB 586
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s6447 => state := s6448;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (635, 12)); -- offset MSB 587
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6448 => state := s6449; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6449 => 			--4
	if (fixed2floatrdy = '1') then state := s6450;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6449; end if;
when s6450 => state := s6451; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6451 => 			--6
	if (mulfprdy = '1') then state := s6452;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6451; end if;
when s6452 => state := s6453; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6453 => 			--8
	if (mulfprdy = '1') then state := s6454;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6453; end if;
when s6454 => state := s6455; 	--9
	mulfpsclr <= '0';
when s6455 => state := s6456; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6456 => 			--11
	if (mulfprdy = '1') then state := s6457;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6456; end if;
when s6457 => state := s6458; 	--12
	mulfpsclr <= '0';
when s6458 => state := s6459; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6459 => 			--14
	if (addfprdy = '1') then state := s6460;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6459; end if;
when s6460 => state := s6461; 	--15
	addfpsclr <= '0';
when s6461 => state := s6462; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6462 => 			--17
	if (addfprdy = '1') then state := s6463;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6462; end if;
when s6463 => state := s6464; 	--18
	addfpsclr <= '0';
when s6464 => state := s6465; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6465 => 			--20
	if (addfprdy = '1') then state := s6466;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6465; end if;
when s6466 => state := s6467; 	--21
	addfpsclr <= '0';
when s6467 => state := s6468; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (349, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6468 => state := s6469; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (636, 12)); -- offset LSB 588
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s6469 => state := s6470;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (637, 12)); -- offset MSB 589
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6470 => state := s6471; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6471 => 			--4
	if (fixed2floatrdy = '1') then state := s6472;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6471; end if;
when s6472 => state := s6473; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6473 => 			--6
	if (mulfprdy = '1') then state := s6474;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6473; end if;
when s6474 => state := s6475; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6475 => 			--8
	if (mulfprdy = '1') then state := s6476;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6475; end if;
when s6476 => state := s6477; 	--9
	mulfpsclr <= '0';
when s6477 => state := s6478; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6478 => 			--11
	if (mulfprdy = '1') then state := s6479;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6478; end if;
when s6479 => state := s6480; 	--12
	mulfpsclr <= '0';
when s6480 => state := s6481; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6481 => 			--14
	if (addfprdy = '1') then state := s6482;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6481; end if;
when s6482 => state := s6483; 	--15
	addfpsclr <= '0';
when s6483 => state := s6484; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6484 => 			--17
	if (addfprdy = '1') then state := s6485;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6484; end if;
when s6485 => state := s6486; 	--18
	addfpsclr <= '0';
when s6486 => state := s6487; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6487 => 			--20
	if (addfprdy = '1') then state := s6488;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6487; end if;
when s6488 => state := s6489; 	--21
	addfpsclr <= '0';
when s6489 => state := s6490; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (350, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6490 => state := s6491; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (638, 12)); -- offset LSB 590
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s6491 => state := s6492;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (639, 12)); -- offset MSB 591
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6492 => state := s6493; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6493 => 			--4
	if (fixed2floatrdy = '1') then state := s6494;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6493; end if;
when s6494 => state := s6495; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6495 => 			--6
	if (mulfprdy = '1') then state := s6496;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6495; end if;
when s6496 => state := s6497; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6497 => 			--8
	if (mulfprdy = '1') then state := s6498;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6497; end if;
when s6498 => state := s6499; 	--9
	mulfpsclr <= '0';
when s6499 => state := s6500; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6500 => 			--11
	if (mulfprdy = '1') then state := s6501;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6500; end if;
when s6501 => state := s6502; 	--12
	mulfpsclr <= '0';
when s6502 => state := s6503; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6503 => 			--14
	if (addfprdy = '1') then state := s6504;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6503; end if;
when s6504 => state := s6505; 	--15
	addfpsclr <= '0';
when s6505 => state := s6506; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6506 => 			--17
	if (addfprdy = '1') then state := s6507;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6506; end if;
when s6507 => state := s6508; 	--18
	addfpsclr <= '0';
when s6508 => state := s6509; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6509 => 			--20
	if (addfprdy = '1') then state := s6510;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6509; end if;
when s6510 => state := s6511; 	--21
	addfpsclr <= '0';
when s6511 => state := s6512; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (351, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6512 => state := s6513; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (640, 12)); -- offset LSB 592
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s6513 => state := s6514;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (641, 12)); -- offset MSB 593
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6514 => state := s6515; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6515 => 			--4
	if (fixed2floatrdy = '1') then state := s6516;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6515; end if;
when s6516 => state := s6517; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6517 => 			--6
	if (mulfprdy = '1') then state := s6518;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6517; end if;
when s6518 => state := s6519; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6519 => 			--8
	if (mulfprdy = '1') then state := s6520;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6519; end if;
when s6520 => state := s6521; 	--9
	mulfpsclr <= '0';
when s6521 => state := s6522; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6522 => 			--11
	if (mulfprdy = '1') then state := s6523;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6522; end if;
when s6523 => state := s6524; 	--12
	mulfpsclr <= '0';
when s6524 => state := s6525; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6525 => 			--14
	if (addfprdy = '1') then state := s6526;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6525; end if;
when s6526 => state := s6527; 	--15
	addfpsclr <= '0';
when s6527 => state := s6528; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6528 => 			--17
	if (addfprdy = '1') then state := s6529;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6528; end if;
when s6529 => state := s6530; 	--18
	addfpsclr <= '0';
when s6530 => state := s6531; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6531 => 			--20
	if (addfprdy = '1') then state := s6532;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6531; end if;
when s6532 => state := s6533; 	--21
	addfpsclr <= '0';
when s6533 => state := s6534; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (352, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6534 => state := s6535; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (642, 12)); -- offset LSB 594
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s6535 => state := s6536;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (643, 12)); -- offset MSB 595
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6536 => state := s6537; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6537 => 			--4
	if (fixed2floatrdy = '1') then state := s6538;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6537; end if;
when s6538 => state := s6539; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6539 => 			--6
	if (mulfprdy = '1') then state := s6540;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6539; end if;
when s6540 => state := s6541; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6541 => 			--8
	if (mulfprdy = '1') then state := s6542;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6541; end if;
when s6542 => state := s6543; 	--9
	mulfpsclr <= '0';
when s6543 => state := s6544; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6544 => 			--11
	if (mulfprdy = '1') then state := s6545;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6544; end if;
when s6545 => state := s6546; 	--12
	mulfpsclr <= '0';
when s6546 => state := s6547; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6547 => 			--14
	if (addfprdy = '1') then state := s6548;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6547; end if;
when s6548 => state := s6549; 	--15
	addfpsclr <= '0';
when s6549 => state := s6550; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6550 => 			--17
	if (addfprdy = '1') then state := s6551;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6550; end if;
when s6551 => state := s6552; 	--18
	addfpsclr <= '0';
when s6552 => state := s6553; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6553 => 			--20
	if (addfprdy = '1') then state := s6554;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6553; end if;
when s6554 => state := s6555; 	--21
	addfpsclr <= '0';
when s6555 => state := s6556; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (353, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6556 => state := s6557; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (644, 12)); -- offset LSB 596
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s6557 => state := s6558;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (645, 12)); -- offset MSB 597
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6558 => state := s6559; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6559 => 			--4
	if (fixed2floatrdy = '1') then state := s6560;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6559; end if;
when s6560 => state := s6561; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6561 => 			--6
	if (mulfprdy = '1') then state := s6562;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6561; end if;
when s6562 => state := s6563; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6563 => 			--8
	if (mulfprdy = '1') then state := s6564;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6563; end if;
when s6564 => state := s6565; 	--9
	mulfpsclr <= '0';
when s6565 => state := s6566; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6566 => 			--11
	if (mulfprdy = '1') then state := s6567;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6566; end if;
when s6567 => state := s6568; 	--12
	mulfpsclr <= '0';
when s6568 => state := s6569; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6569 => 			--14
	if (addfprdy = '1') then state := s6570;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6569; end if;
when s6570 => state := s6571; 	--15
	addfpsclr <= '0';
when s6571 => state := s6572; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6572 => 			--17
	if (addfprdy = '1') then state := s6573;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6572; end if;
when s6573 => state := s6574; 	--18
	addfpsclr <= '0';
when s6574 => state := s6575; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6575 => 			--20
	if (addfprdy = '1') then state := s6576;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6575; end if;
when s6576 => state := s6577; 	--21
	addfpsclr <= '0';
when s6577 => state := s6578; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (354, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6578 => state := s6579; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (646, 12)); -- offset LSB 598
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s6579 => state := s6580;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (647, 12)); -- offset MSB 599
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6580 => state := s6581; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6581 => 			--4
	if (fixed2floatrdy = '1') then state := s6582;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6581; end if;
when s6582 => state := s6583; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6583 => 			--6
	if (mulfprdy = '1') then state := s6584;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6583; end if;
when s6584 => state := s6585; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6585 => 			--8
	if (mulfprdy = '1') then state := s6586;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6585; end if;
when s6586 => state := s6587; 	--9
	mulfpsclr <= '0';
when s6587 => state := s6588; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6588 => 			--11
	if (mulfprdy = '1') then state := s6589;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6588; end if;
when s6589 => state := s6590; 	--12
	mulfpsclr <= '0';
when s6590 => state := s6591; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6591 => 			--14
	if (addfprdy = '1') then state := s6592;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6591; end if;
when s6592 => state := s6593; 	--15
	addfpsclr <= '0';
when s6593 => state := s6594; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6594 => 			--17
	if (addfprdy = '1') then state := s6595;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6594; end if;
when s6595 => state := s6596; 	--18
	addfpsclr <= '0';
when s6596 => state := s6597; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6597 => 			--20
	if (addfprdy = '1') then state := s6598;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6597; end if;
when s6598 => state := s6599; 	--21
	addfpsclr <= '0';
when s6599 => state := s6600; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (355, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6600 => state := s6601; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (648, 12)); -- offset LSB 600
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s6601 => state := s6602;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (649, 12)); -- offset MSB 601
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6602 => state := s6603; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6603 => 			--4
	if (fixed2floatrdy = '1') then state := s6604;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6603; end if;
when s6604 => state := s6605; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6605 => 			--6
	if (mulfprdy = '1') then state := s6606;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6605; end if;
when s6606 => state := s6607; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6607 => 			--8
	if (mulfprdy = '1') then state := s6608;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6607; end if;
when s6608 => state := s6609; 	--9
	mulfpsclr <= '0';
when s6609 => state := s6610; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6610 => 			--11
	if (mulfprdy = '1') then state := s6611;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6610; end if;
when s6611 => state := s6612; 	--12
	mulfpsclr <= '0';
when s6612 => state := s6613; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6613 => 			--14
	if (addfprdy = '1') then state := s6614;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6613; end if;
when s6614 => state := s6615; 	--15
	addfpsclr <= '0';
when s6615 => state := s6616; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6616 => 			--17
	if (addfprdy = '1') then state := s6617;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6616; end if;
when s6617 => state := s6618; 	--18
	addfpsclr <= '0';
when s6618 => state := s6619; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6619 => 			--20
	if (addfprdy = '1') then state := s6620;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6619; end if;
when s6620 => state := s6621; 	--21
	addfpsclr <= '0';
when s6621 => state := s6622; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (356, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6622 => state := s6623; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (650, 12)); -- offset LSB 602
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s6623 => state := s6624;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (651, 12)); -- offset MSB 603
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6624 => state := s6625; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6625 => 			--4
	if (fixed2floatrdy = '1') then state := s6626;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6625; end if;
when s6626 => state := s6627; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6627 => 			--6
	if (mulfprdy = '1') then state := s6628;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6627; end if;
when s6628 => state := s6629; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6629 => 			--8
	if (mulfprdy = '1') then state := s6630;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6629; end if;
when s6630 => state := s6631; 	--9
	mulfpsclr <= '0';
when s6631 => state := s6632; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6632 => 			--11
	if (mulfprdy = '1') then state := s6633;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6632; end if;
when s6633 => state := s6634; 	--12
	mulfpsclr <= '0';
when s6634 => state := s6635; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6635 => 			--14
	if (addfprdy = '1') then state := s6636;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6635; end if;
when s6636 => state := s6637; 	--15
	addfpsclr <= '0';
when s6637 => state := s6638; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6638 => 			--17
	if (addfprdy = '1') then state := s6639;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6638; end if;
when s6639 => state := s6640; 	--18
	addfpsclr <= '0';
when s6640 => state := s6641; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6641 => 			--20
	if (addfprdy = '1') then state := s6642;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6641; end if;
when s6642 => state := s6643; 	--21
	addfpsclr <= '0';
when s6643 => state := s6644; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (357, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6644 => state := s6645; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (652, 12)); -- offset LSB 604
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s6645 => state := s6646;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (653, 12)); -- offset MSB 605
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6646 => state := s6647; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6647 => 			--4
	if (fixed2floatrdy = '1') then state := s6648;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6647; end if;
when s6648 => state := s6649; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6649 => 			--6
	if (mulfprdy = '1') then state := s6650;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6649; end if;
when s6650 => state := s6651; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6651 => 			--8
	if (mulfprdy = '1') then state := s6652;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6651; end if;
when s6652 => state := s6653; 	--9
	mulfpsclr <= '0';
when s6653 => state := s6654; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6654 => 			--11
	if (mulfprdy = '1') then state := s6655;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6654; end if;
when s6655 => state := s6656; 	--12
	mulfpsclr <= '0';
when s6656 => state := s6657; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6657 => 			--14
	if (addfprdy = '1') then state := s6658;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6657; end if;
when s6658 => state := s6659; 	--15
	addfpsclr <= '0';
when s6659 => state := s6660; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6660 => 			--17
	if (addfprdy = '1') then state := s6661;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6660; end if;
when s6661 => state := s6662; 	--18
	addfpsclr <= '0';
when s6662 => state := s6663; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6663 => 			--20
	if (addfprdy = '1') then state := s6664;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6663; end if;
when s6664 => state := s6665; 	--21
	addfpsclr <= '0';
when s6665 => state := s6666; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (358, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6666 => state := s6667; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (654, 12)); -- offset LSB 606
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s6667 => state := s6668;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (655, 12)); -- offset MSB 607
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6668 => state := s6669; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6669 => 			--4
	if (fixed2floatrdy = '1') then state := s6670;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6669; end if;
when s6670 => state := s6671; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6671 => 			--6
	if (mulfprdy = '1') then state := s6672;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6671; end if;
when s6672 => state := s6673; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6673 => 			--8
	if (mulfprdy = '1') then state := s6674;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6673; end if;
when s6674 => state := s6675; 	--9
	mulfpsclr <= '0';
when s6675 => state := s6676; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6676 => 			--11
	if (mulfprdy = '1') then state := s6677;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6676; end if;
when s6677 => state := s6678; 	--12
	mulfpsclr <= '0';
when s6678 => state := s6679; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6679 => 			--14
	if (addfprdy = '1') then state := s6680;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6679; end if;
when s6680 => state := s6681; 	--15
	addfpsclr <= '0';
when s6681 => state := s6682; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6682 => 			--17
	if (addfprdy = '1') then state := s6683;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6682; end if;
when s6683 => state := s6684; 	--18
	addfpsclr <= '0';
when s6684 => state := s6685; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6685 => 			--20
	if (addfprdy = '1') then state := s6686;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6685; end if;
when s6686 => state := s6687; 	--21
	addfpsclr <= '0';
when s6687 => state := s6688; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (359, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6688 => state := s6689; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (656, 12)); -- offset LSB 608
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s6689 => state := s6690;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (657, 12)); -- offset MSB 609
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6690 => state := s6691; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6691 => 			--4
	if (fixed2floatrdy = '1') then state := s6692;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6691; end if;
when s6692 => state := s6693; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6693 => 			--6
	if (mulfprdy = '1') then state := s6694;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6693; end if;
when s6694 => state := s6695; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6695 => 			--8
	if (mulfprdy = '1') then state := s6696;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6695; end if;
when s6696 => state := s6697; 	--9
	mulfpsclr <= '0';
when s6697 => state := s6698; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6698 => 			--11
	if (mulfprdy = '1') then state := s6699;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6698; end if;
when s6699 => state := s6700; 	--12
	mulfpsclr <= '0';
when s6700 => state := s6701; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6701 => 			--14
	if (addfprdy = '1') then state := s6702;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6701; end if;
when s6702 => state := s6703; 	--15
	addfpsclr <= '0';
when s6703 => state := s6704; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6704 => 			--17
	if (addfprdy = '1') then state := s6705;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6704; end if;
when s6705 => state := s6706; 	--18
	addfpsclr <= '0';
when s6706 => state := s6707; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6707 => 			--20
	if (addfprdy = '1') then state := s6708;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6707; end if;
when s6708 => state := s6709; 	--21
	addfpsclr <= '0';
when s6709 => state := s6710; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (360, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6710 => state := s6711; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (658, 12)); -- offset LSB 610
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s6711 => state := s6712;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (659, 12)); -- offset MSB 611
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6712 => state := s6713; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6713 => 			--4
	if (fixed2floatrdy = '1') then state := s6714;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6713; end if;
when s6714 => state := s6715; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6715 => 			--6
	if (mulfprdy = '1') then state := s6716;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6715; end if;
when s6716 => state := s6717; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6717 => 			--8
	if (mulfprdy = '1') then state := s6718;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6717; end if;
when s6718 => state := s6719; 	--9
	mulfpsclr <= '0';
when s6719 => state := s6720; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6720 => 			--11
	if (mulfprdy = '1') then state := s6721;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6720; end if;
when s6721 => state := s6722; 	--12
	mulfpsclr <= '0';
when s6722 => state := s6723; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6723 => 			--14
	if (addfprdy = '1') then state := s6724;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6723; end if;
when s6724 => state := s6725; 	--15
	addfpsclr <= '0';
when s6725 => state := s6726; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6726 => 			--17
	if (addfprdy = '1') then state := s6727;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6726; end if;
when s6727 => state := s6728; 	--18
	addfpsclr <= '0';
when s6728 => state := s6729; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6729 => 			--20
	if (addfprdy = '1') then state := s6730;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6729; end if;
when s6730 => state := s6731; 	--21
	addfpsclr <= '0';
when s6731 => state := s6732; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (361, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6732 => state := s6733; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (660, 12)); -- offset LSB 612
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s6733 => state := s6734;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (661, 12)); -- offset MSB 613
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6734 => state := s6735; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6735 => 			--4
	if (fixed2floatrdy = '1') then state := s6736;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6735; end if;
when s6736 => state := s6737; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6737 => 			--6
	if (mulfprdy = '1') then state := s6738;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6737; end if;
when s6738 => state := s6739; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6739 => 			--8
	if (mulfprdy = '1') then state := s6740;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6739; end if;
when s6740 => state := s6741; 	--9
	mulfpsclr <= '0';
when s6741 => state := s6742; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6742 => 			--11
	if (mulfprdy = '1') then state := s6743;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6742; end if;
when s6743 => state := s6744; 	--12
	mulfpsclr <= '0';
when s6744 => state := s6745; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6745 => 			--14
	if (addfprdy = '1') then state := s6746;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6745; end if;
when s6746 => state := s6747; 	--15
	addfpsclr <= '0';
when s6747 => state := s6748; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6748 => 			--17
	if (addfprdy = '1') then state := s6749;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6748; end if;
when s6749 => state := s6750; 	--18
	addfpsclr <= '0';
when s6750 => state := s6751; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6751 => 			--20
	if (addfprdy = '1') then state := s6752;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6751; end if;
when s6752 => state := s6753; 	--21
	addfpsclr <= '0';
when s6753 => state := s6754; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (362, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6754 => state := s6755; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (662, 12)); -- offset LSB 614
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s6755 => state := s6756;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (663, 12)); -- offset MSB 615
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6756 => state := s6757; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6757 => 			--4
	if (fixed2floatrdy = '1') then state := s6758;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6757; end if;
when s6758 => state := s6759; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6759 => 			--6
	if (mulfprdy = '1') then state := s6760;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6759; end if;
when s6760 => state := s6761; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6761 => 			--8
	if (mulfprdy = '1') then state := s6762;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6761; end if;
when s6762 => state := s6763; 	--9
	mulfpsclr <= '0';
when s6763 => state := s6764; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6764 => 			--11
	if (mulfprdy = '1') then state := s6765;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6764; end if;
when s6765 => state := s6766; 	--12
	mulfpsclr <= '0';
when s6766 => state := s6767; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6767 => 			--14
	if (addfprdy = '1') then state := s6768;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6767; end if;
when s6768 => state := s6769; 	--15
	addfpsclr <= '0';
when s6769 => state := s6770; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6770 => 			--17
	if (addfprdy = '1') then state := s6771;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6770; end if;
when s6771 => state := s6772; 	--18
	addfpsclr <= '0';
when s6772 => state := s6773; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6773 => 			--20
	if (addfprdy = '1') then state := s6774;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6773; end if;
when s6774 => state := s6775; 	--21
	addfpsclr <= '0';
when s6775 => state := s6776; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (363, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6776 => state := s6777; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (664, 12)); -- offset LSB 616
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s6777 => state := s6778;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (665, 12)); -- offset MSB 617
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6778 => state := s6779; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6779 => 			--4
	if (fixed2floatrdy = '1') then state := s6780;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6779; end if;
when s6780 => state := s6781; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6781 => 			--6
	if (mulfprdy = '1') then state := s6782;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6781; end if;
when s6782 => state := s6783; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6783 => 			--8
	if (mulfprdy = '1') then state := s6784;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6783; end if;
when s6784 => state := s6785; 	--9
	mulfpsclr <= '0';
when s6785 => state := s6786; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6786 => 			--11
	if (mulfprdy = '1') then state := s6787;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6786; end if;
when s6787 => state := s6788; 	--12
	mulfpsclr <= '0';
when s6788 => state := s6789; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6789 => 			--14
	if (addfprdy = '1') then state := s6790;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6789; end if;
when s6790 => state := s6791; 	--15
	addfpsclr <= '0';
when s6791 => state := s6792; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6792 => 			--17
	if (addfprdy = '1') then state := s6793;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6792; end if;
when s6793 => state := s6794; 	--18
	addfpsclr <= '0';
when s6794 => state := s6795; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6795 => 			--20
	if (addfprdy = '1') then state := s6796;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6795; end if;
when s6796 => state := s6797; 	--21
	addfpsclr <= '0';
when s6797 => state := s6798; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (364, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6798 => state := s6799; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (666, 12)); -- offset LSB 618
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s6799 => state := s6800;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (667, 12)); -- offset MSB 619
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6800 => state := s6801; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6801 => 			--4
	if (fixed2floatrdy = '1') then state := s6802;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6801; end if;
when s6802 => state := s6803; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6803 => 			--6
	if (mulfprdy = '1') then state := s6804;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6803; end if;
when s6804 => state := s6805; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6805 => 			--8
	if (mulfprdy = '1') then state := s6806;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6805; end if;
when s6806 => state := s6807; 	--9
	mulfpsclr <= '0';
when s6807 => state := s6808; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6808 => 			--11
	if (mulfprdy = '1') then state := s6809;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6808; end if;
when s6809 => state := s6810; 	--12
	mulfpsclr <= '0';
when s6810 => state := s6811; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6811 => 			--14
	if (addfprdy = '1') then state := s6812;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6811; end if;
when s6812 => state := s6813; 	--15
	addfpsclr <= '0';
when s6813 => state := s6814; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6814 => 			--17
	if (addfprdy = '1') then state := s6815;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6814; end if;
when s6815 => state := s6816; 	--18
	addfpsclr <= '0';
when s6816 => state := s6817; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6817 => 			--20
	if (addfprdy = '1') then state := s6818;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6817; end if;
when s6818 => state := s6819; 	--21
	addfpsclr <= '0';
when s6819 => state := s6820; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (365, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6820 => state := s6821; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (668, 12)); -- offset LSB 620
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s6821 => state := s6822;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (669, 12)); -- offset MSB 621
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6822 => state := s6823; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6823 => 			--4
	if (fixed2floatrdy = '1') then state := s6824;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6823; end if;
when s6824 => state := s6825; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6825 => 			--6
	if (mulfprdy = '1') then state := s6826;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6825; end if;
when s6826 => state := s6827; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6827 => 			--8
	if (mulfprdy = '1') then state := s6828;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6827; end if;
when s6828 => state := s6829; 	--9
	mulfpsclr <= '0';
when s6829 => state := s6830; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6830 => 			--11
	if (mulfprdy = '1') then state := s6831;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6830; end if;
when s6831 => state := s6832; 	--12
	mulfpsclr <= '0';
when s6832 => state := s6833; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6833 => 			--14
	if (addfprdy = '1') then state := s6834;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6833; end if;
when s6834 => state := s6835; 	--15
	addfpsclr <= '0';
when s6835 => state := s6836; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6836 => 			--17
	if (addfprdy = '1') then state := s6837;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6836; end if;
when s6837 => state := s6838; 	--18
	addfpsclr <= '0';
when s6838 => state := s6839; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6839 => 			--20
	if (addfprdy = '1') then state := s6840;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6839; end if;
when s6840 => state := s6841; 	--21
	addfpsclr <= '0';
when s6841 => state := s6842; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (366, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6842 => state := s6843; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (670, 12)); -- offset LSB 622
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s6843 => state := s6844;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (671, 12)); -- offset MSB 623
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6844 => state := s6845; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6845 => 			--4
	if (fixed2floatrdy = '1') then state := s6846;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6845; end if;
when s6846 => state := s6847; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6847 => 			--6
	if (mulfprdy = '1') then state := s6848;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6847; end if;
when s6848 => state := s6849; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6849 => 			--8
	if (mulfprdy = '1') then state := s6850;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6849; end if;
when s6850 => state := s6851; 	--9
	mulfpsclr <= '0';
when s6851 => state := s6852; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6852 => 			--11
	if (mulfprdy = '1') then state := s6853;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6852; end if;
when s6853 => state := s6854; 	--12
	mulfpsclr <= '0';
when s6854 => state := s6855; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6855 => 			--14
	if (addfprdy = '1') then state := s6856;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6855; end if;
when s6856 => state := s6857; 	--15
	addfpsclr <= '0';
when s6857 => state := s6858; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6858 => 			--17
	if (addfprdy = '1') then state := s6859;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6858; end if;
when s6859 => state := s6860; 	--18
	addfpsclr <= '0';
when s6860 => state := s6861; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6861 => 			--20
	if (addfprdy = '1') then state := s6862;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6861; end if;
when s6862 => state := s6863; 	--21
	addfpsclr <= '0';
when s6863 => state := s6864; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (367, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6864 => state := s6865; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (672, 12)); -- offset LSB 624
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s6865 => state := s6866;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (673, 12)); -- offset MSB 625
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6866 => state := s6867; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6867 => 			--4
	if (fixed2floatrdy = '1') then state := s6868;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6867; end if;
when s6868 => state := s6869; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6869 => 			--6
	if (mulfprdy = '1') then state := s6870;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6869; end if;
when s6870 => state := s6871; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6871 => 			--8
	if (mulfprdy = '1') then state := s6872;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6871; end if;
when s6872 => state := s6873; 	--9
	mulfpsclr <= '0';
when s6873 => state := s6874; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6874 => 			--11
	if (mulfprdy = '1') then state := s6875;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6874; end if;
when s6875 => state := s6876; 	--12
	mulfpsclr <= '0';
when s6876 => state := s6877; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6877 => 			--14
	if (addfprdy = '1') then state := s6878;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6877; end if;
when s6878 => state := s6879; 	--15
	addfpsclr <= '0';
when s6879 => state := s6880; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6880 => 			--17
	if (addfprdy = '1') then state := s6881;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6880; end if;
when s6881 => state := s6882; 	--18
	addfpsclr <= '0';
when s6882 => state := s6883; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6883 => 			--20
	if (addfprdy = '1') then state := s6884;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6883; end if;
when s6884 => state := s6885; 	--21
	addfpsclr <= '0';
when s6885 => state := s6886; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (368, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6886 => state := s6887; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (674, 12)); -- offset LSB 626
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s6887 => state := s6888;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (675, 12)); -- offset MSB 627
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6888 => state := s6889; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6889 => 			--4
	if (fixed2floatrdy = '1') then state := s6890;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6889; end if;
when s6890 => state := s6891; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6891 => 			--6
	if (mulfprdy = '1') then state := s6892;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6891; end if;
when s6892 => state := s6893; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6893 => 			--8
	if (mulfprdy = '1') then state := s6894;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6893; end if;
when s6894 => state := s6895; 	--9
	mulfpsclr <= '0';
when s6895 => state := s6896; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6896 => 			--11
	if (mulfprdy = '1') then state := s6897;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6896; end if;
when s6897 => state := s6898; 	--12
	mulfpsclr <= '0';
when s6898 => state := s6899; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6899 => 			--14
	if (addfprdy = '1') then state := s6900;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6899; end if;
when s6900 => state := s6901; 	--15
	addfpsclr <= '0';
when s6901 => state := s6902; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6902 => 			--17
	if (addfprdy = '1') then state := s6903;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6902; end if;
when s6903 => state := s6904; 	--18
	addfpsclr <= '0';
when s6904 => state := s6905; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6905 => 			--20
	if (addfprdy = '1') then state := s6906;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6905; end if;
when s6906 => state := s6907; 	--21
	addfpsclr <= '0';
when s6907 => state := s6908; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (369, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6908 => state := s6909; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (676, 12)); -- offset LSB 628
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s6909 => state := s6910;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (677, 12)); -- offset MSB 629
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6910 => state := s6911; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6911 => 			--4
	if (fixed2floatrdy = '1') then state := s6912;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6911; end if;
when s6912 => state := s6913; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6913 => 			--6
	if (mulfprdy = '1') then state := s6914;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6913; end if;
when s6914 => state := s6915; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6915 => 			--8
	if (mulfprdy = '1') then state := s6916;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6915; end if;
when s6916 => state := s6917; 	--9
	mulfpsclr <= '0';
when s6917 => state := s6918; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6918 => 			--11
	if (mulfprdy = '1') then state := s6919;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6918; end if;
when s6919 => state := s6920; 	--12
	mulfpsclr <= '0';
when s6920 => state := s6921; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6921 => 			--14
	if (addfprdy = '1') then state := s6922;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6921; end if;
when s6922 => state := s6923; 	--15
	addfpsclr <= '0';
when s6923 => state := s6924; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6924 => 			--17
	if (addfprdy = '1') then state := s6925;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6924; end if;
when s6925 => state := s6926; 	--18
	addfpsclr <= '0';
when s6926 => state := s6927; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6927 => 			--20
	if (addfprdy = '1') then state := s6928;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6927; end if;
when s6928 => state := s6929; 	--21
	addfpsclr <= '0';
when s6929 => state := s6930; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (370, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6930 => state := s6931; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (678, 12)); -- offset LSB 630
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s6931 => state := s6932;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (679, 12)); -- offset MSB 631
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6932 => state := s6933; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6933 => 			--4
	if (fixed2floatrdy = '1') then state := s6934;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6933; end if;
when s6934 => state := s6935; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6935 => 			--6
	if (mulfprdy = '1') then state := s6936;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6935; end if;
when s6936 => state := s6937; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6937 => 			--8
	if (mulfprdy = '1') then state := s6938;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6937; end if;
when s6938 => state := s6939; 	--9
	mulfpsclr <= '0';
when s6939 => state := s6940; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6940 => 			--11
	if (mulfprdy = '1') then state := s6941;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6940; end if;
when s6941 => state := s6942; 	--12
	mulfpsclr <= '0';
when s6942 => state := s6943; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6943 => 			--14
	if (addfprdy = '1') then state := s6944;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6943; end if;
when s6944 => state := s6945; 	--15
	addfpsclr <= '0';
when s6945 => state := s6946; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6946 => 			--17
	if (addfprdy = '1') then state := s6947;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6946; end if;
when s6947 => state := s6948; 	--18
	addfpsclr <= '0';
when s6948 => state := s6949; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6949 => 			--20
	if (addfprdy = '1') then state := s6950;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6949; end if;
when s6950 => state := s6951; 	--21
	addfpsclr <= '0';
when s6951 => state := s6952; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (371, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6952 => state := s6953; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (680, 12)); -- offset LSB 632
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s6953 => state := s6954;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (681, 12)); -- offset MSB 633
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6954 => state := s6955; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6955 => 			--4
	if (fixed2floatrdy = '1') then state := s6956;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6955; end if;
when s6956 => state := s6957; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6957 => 			--6
	if (mulfprdy = '1') then state := s6958;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6957; end if;
when s6958 => state := s6959; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6959 => 			--8
	if (mulfprdy = '1') then state := s6960;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6959; end if;
when s6960 => state := s6961; 	--9
	mulfpsclr <= '0';
when s6961 => state := s6962; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6962 => 			--11
	if (mulfprdy = '1') then state := s6963;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6962; end if;
when s6963 => state := s6964; 	--12
	mulfpsclr <= '0';
when s6964 => state := s6965; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6965 => 			--14
	if (addfprdy = '1') then state := s6966;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6965; end if;
when s6966 => state := s6967; 	--15
	addfpsclr <= '0';
when s6967 => state := s6968; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6968 => 			--17
	if (addfprdy = '1') then state := s6969;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6968; end if;
when s6969 => state := s6970; 	--18
	addfpsclr <= '0';
when s6970 => state := s6971; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6971 => 			--20
	if (addfprdy = '1') then state := s6972;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6971; end if;
when s6972 => state := s6973; 	--21
	addfpsclr <= '0';
when s6973 => state := s6974; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (372, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6974 => state := s6975; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (682, 12)); -- offset LSB 634
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s6975 => state := s6976;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (683, 12)); -- offset MSB 635
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6976 => state := s6977; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6977 => 			--4
	if (fixed2floatrdy = '1') then state := s6978;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6977; end if;
when s6978 => state := s6979; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s6979 => 			--6
	if (mulfprdy = '1') then state := s6980;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6979; end if;
when s6980 => state := s6981; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s6981 => 			--8
	if (mulfprdy = '1') then state := s6982;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6981; end if;
when s6982 => state := s6983; 	--9
	mulfpsclr <= '0';
when s6983 => state := s6984; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s6984 => 			--11
	if (mulfprdy = '1') then state := s6985;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s6984; end if;
when s6985 => state := s6986; 	--12
	mulfpsclr <= '0';
when s6986 => state := s6987; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s6987 => 			--14
	if (addfprdy = '1') then state := s6988;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6987; end if;
when s6988 => state := s6989; 	--15
	addfpsclr <= '0';
when s6989 => state := s6990; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s6990 => 			--17
	if (addfprdy = '1') then state := s6991;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6990; end if;
when s6991 => state := s6992; 	--18
	addfpsclr <= '0';
when s6992 => state := s6993; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s6993 => 			--20
	if (addfprdy = '1') then state := s6994;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s6993; end if;
when s6994 => state := s6995; 	--21
	addfpsclr <= '0';
when s6995 => state := s6996; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (373, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s6996 => state := s6997; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (684, 12)); -- offset LSB 636
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s6997 => state := s6998;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (685, 12)); -- offset MSB 637
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s6998 => state := s6999; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s6999 => 			--4
	if (fixed2floatrdy = '1') then state := s7000;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s6999; end if;
when s7000 => state := s7001; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7001 => 			--6
	if (mulfprdy = '1') then state := s7002;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7001; end if;
when s7002 => state := s7003; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7003 => 			--8
	if (mulfprdy = '1') then state := s7004;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7003; end if;
when s7004 => state := s7005; 	--9
	mulfpsclr <= '0';
when s7005 => state := s7006; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7006 => 			--11
	if (mulfprdy = '1') then state := s7007;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7006; end if;
when s7007 => state := s7008; 	--12
	mulfpsclr <= '0';
when s7008 => state := s7009; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7009 => 			--14
	if (addfprdy = '1') then state := s7010;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7009; end if;
when s7010 => state := s7011; 	--15
	addfpsclr <= '0';
when s7011 => state := s7012; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7012 => 			--17
	if (addfprdy = '1') then state := s7013;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7012; end if;
when s7013 => state := s7014; 	--18
	addfpsclr <= '0';
when s7014 => state := s7015; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7015 => 			--20
	if (addfprdy = '1') then state := s7016;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7015; end if;
when s7016 => state := s7017; 	--21
	addfpsclr <= '0';
when s7017 => state := s7018; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (374, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7018 => state := s7019; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (686, 12)); -- offset LSB 638
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s7019 => state := s7020;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (687, 12)); -- offset MSB 639
	addra <= std_logic_vector (to_unsigned (9, 10)); -- OCCrowI 9
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7020 => state := s7021; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7021 => 			--4
	if (fixed2floatrdy = '1') then state := s7022;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7021; end if;
when s7022 => state := s7023; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7023 => 			--6
	if (mulfprdy = '1') then state := s7024;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7023; end if;
when s7024 => state := s7025; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7025 => 			--8
	if (mulfprdy = '1') then state := s7026;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7025; end if;
when s7026 => state := s7027; 	--9
	mulfpsclr <= '0';
when s7027 => state := s7028; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7028 => 			--11
	if (mulfprdy = '1') then state := s7029;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7028; end if;
when s7029 => state := s7030; 	--12
	mulfpsclr <= '0';
when s7030 => state := s7031; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7031 => 			--14
	if (addfprdy = '1') then state := s7032;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7031; end if;
when s7032 => state := s7033; 	--15
	addfpsclr <= '0';
when s7033 => state := s7034; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7034 => 			--17
	if (addfprdy = '1') then state := s7035;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7034; end if;
when s7035 => state := s7036; 	--18
	addfpsclr <= '0';
when s7036 => state := s7037; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7037 => 			--20
	if (addfprdy = '1') then state := s7038;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7037; end if;
when s7038 => state := s7039; 	--21
	addfpsclr <= '0';
when s7039 => state := s7040; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (375, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7040 => state := s7041; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (688, 12)); -- offset LSB 640
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s7041 => state := s7042;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (689, 12)); -- offset MSB 641
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7042 => state := s7043; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7043 => 			--4
	if (fixed2floatrdy = '1') then state := s7044;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7043; end if;
when s7044 => state := s7045; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7045 => 			--6
	if (mulfprdy = '1') then state := s7046;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7045; end if;
when s7046 => state := s7047; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7047 => 			--8
	if (mulfprdy = '1') then state := s7048;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7047; end if;
when s7048 => state := s7049; 	--9
	mulfpsclr <= '0';
when s7049 => state := s7050; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7050 => 			--11
	if (mulfprdy = '1') then state := s7051;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7050; end if;
when s7051 => state := s7052; 	--12
	mulfpsclr <= '0';
when s7052 => state := s7053; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7053 => 			--14
	if (addfprdy = '1') then state := s7054;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7053; end if;
when s7054 => state := s7055; 	--15
	addfpsclr <= '0';
when s7055 => state := s7056; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7056 => 			--17
	if (addfprdy = '1') then state := s7057;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7056; end if;
when s7057 => state := s7058; 	--18
	addfpsclr <= '0';
when s7058 => state := s7059; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7059 => 			--20
	if (addfprdy = '1') then state := s7060;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7059; end if;
when s7060 => state := s7061; 	--21
	addfpsclr <= '0';
when s7061 => state := s7062; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (376, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7062 => state := s7063; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (690, 12)); -- offset LSB 642
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s7063 => state := s7064;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (691, 12)); -- offset MSB 643
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7064 => state := s7065; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7065 => 			--4
	if (fixed2floatrdy = '1') then state := s7066;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7065; end if;
when s7066 => state := s7067; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7067 => 			--6
	if (mulfprdy = '1') then state := s7068;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7067; end if;
when s7068 => state := s7069; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7069 => 			--8
	if (mulfprdy = '1') then state := s7070;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7069; end if;
when s7070 => state := s7071; 	--9
	mulfpsclr <= '0';
when s7071 => state := s7072; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7072 => 			--11
	if (mulfprdy = '1') then state := s7073;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7072; end if;
when s7073 => state := s7074; 	--12
	mulfpsclr <= '0';
when s7074 => state := s7075; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7075 => 			--14
	if (addfprdy = '1') then state := s7076;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7075; end if;
when s7076 => state := s7077; 	--15
	addfpsclr <= '0';
when s7077 => state := s7078; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7078 => 			--17
	if (addfprdy = '1') then state := s7079;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7078; end if;
when s7079 => state := s7080; 	--18
	addfpsclr <= '0';
when s7080 => state := s7081; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7081 => 			--20
	if (addfprdy = '1') then state := s7082;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7081; end if;
when s7082 => state := s7083; 	--21
	addfpsclr <= '0';
when s7083 => state := s7084; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (377, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7084 => state := s7085; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (692, 12)); -- offset LSB 644
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s7085 => state := s7086;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (693, 12)); -- offset MSB 645
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7086 => state := s7087; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7087 => 			--4
	if (fixed2floatrdy = '1') then state := s7088;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7087; end if;
when s7088 => state := s7089; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7089 => 			--6
	if (mulfprdy = '1') then state := s7090;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7089; end if;
when s7090 => state := s7091; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7091 => 			--8
	if (mulfprdy = '1') then state := s7092;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7091; end if;
when s7092 => state := s7093; 	--9
	mulfpsclr <= '0';
when s7093 => state := s7094; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7094 => 			--11
	if (mulfprdy = '1') then state := s7095;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7094; end if;
when s7095 => state := s7096; 	--12
	mulfpsclr <= '0';
when s7096 => state := s7097; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7097 => 			--14
	if (addfprdy = '1') then state := s7098;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7097; end if;
when s7098 => state := s7099; 	--15
	addfpsclr <= '0';
when s7099 => state := s7100; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7100 => 			--17
	if (addfprdy = '1') then state := s7101;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7100; end if;
when s7101 => state := s7102; 	--18
	addfpsclr <= '0';
when s7102 => state := s7103; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7103 => 			--20
	if (addfprdy = '1') then state := s7104;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7103; end if;
when s7104 => state := s7105; 	--21
	addfpsclr <= '0';
when s7105 => state := s7106; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (378, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7106 => state := s7107; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (694, 12)); -- offset LSB 646
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s7107 => state := s7108;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (695, 12)); -- offset MSB 647
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7108 => state := s7109; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7109 => 			--4
	if (fixed2floatrdy = '1') then state := s7110;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7109; end if;
when s7110 => state := s7111; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7111 => 			--6
	if (mulfprdy = '1') then state := s7112;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7111; end if;
when s7112 => state := s7113; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7113 => 			--8
	if (mulfprdy = '1') then state := s7114;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7113; end if;
when s7114 => state := s7115; 	--9
	mulfpsclr <= '0';
when s7115 => state := s7116; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7116 => 			--11
	if (mulfprdy = '1') then state := s7117;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7116; end if;
when s7117 => state := s7118; 	--12
	mulfpsclr <= '0';
when s7118 => state := s7119; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7119 => 			--14
	if (addfprdy = '1') then state := s7120;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7119; end if;
when s7120 => state := s7121; 	--15
	addfpsclr <= '0';
when s7121 => state := s7122; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7122 => 			--17
	if (addfprdy = '1') then state := s7123;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7122; end if;
when s7123 => state := s7124; 	--18
	addfpsclr <= '0';
when s7124 => state := s7125; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7125 => 			--20
	if (addfprdy = '1') then state := s7126;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7125; end if;
when s7126 => state := s7127; 	--21
	addfpsclr <= '0';
when s7127 => state := s7128; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (379, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7128 => state := s7129; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (696, 12)); -- offset LSB 648
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s7129 => state := s7130;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (697, 12)); -- offset MSB 649
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7130 => state := s7131; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7131 => 			--4
	if (fixed2floatrdy = '1') then state := s7132;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7131; end if;
when s7132 => state := s7133; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7133 => 			--6
	if (mulfprdy = '1') then state := s7134;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7133; end if;
when s7134 => state := s7135; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7135 => 			--8
	if (mulfprdy = '1') then state := s7136;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7135; end if;
when s7136 => state := s7137; 	--9
	mulfpsclr <= '0';
when s7137 => state := s7138; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7138 => 			--11
	if (mulfprdy = '1') then state := s7139;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7138; end if;
when s7139 => state := s7140; 	--12
	mulfpsclr <= '0';
when s7140 => state := s7141; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7141 => 			--14
	if (addfprdy = '1') then state := s7142;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7141; end if;
when s7142 => state := s7143; 	--15
	addfpsclr <= '0';
when s7143 => state := s7144; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7144 => 			--17
	if (addfprdy = '1') then state := s7145;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7144; end if;
when s7145 => state := s7146; 	--18
	addfpsclr <= '0';
when s7146 => state := s7147; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7147 => 			--20
	if (addfprdy = '1') then state := s7148;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7147; end if;
when s7148 => state := s7149; 	--21
	addfpsclr <= '0';
when s7149 => state := s7150; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (380, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7150 => state := s7151; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (698, 12)); -- offset LSB 650
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s7151 => state := s7152;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (699, 12)); -- offset MSB 651
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7152 => state := s7153; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7153 => 			--4
	if (fixed2floatrdy = '1') then state := s7154;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7153; end if;
when s7154 => state := s7155; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7155 => 			--6
	if (mulfprdy = '1') then state := s7156;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7155; end if;
when s7156 => state := s7157; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7157 => 			--8
	if (mulfprdy = '1') then state := s7158;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7157; end if;
when s7158 => state := s7159; 	--9
	mulfpsclr <= '0';
when s7159 => state := s7160; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7160 => 			--11
	if (mulfprdy = '1') then state := s7161;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7160; end if;
when s7161 => state := s7162; 	--12
	mulfpsclr <= '0';
when s7162 => state := s7163; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7163 => 			--14
	if (addfprdy = '1') then state := s7164;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7163; end if;
when s7164 => state := s7165; 	--15
	addfpsclr <= '0';
when s7165 => state := s7166; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7166 => 			--17
	if (addfprdy = '1') then state := s7167;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7166; end if;
when s7167 => state := s7168; 	--18
	addfpsclr <= '0';
when s7168 => state := s7169; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7169 => 			--20
	if (addfprdy = '1') then state := s7170;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7169; end if;
when s7170 => state := s7171; 	--21
	addfpsclr <= '0';
when s7171 => state := s7172; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (381, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7172 => state := s7173; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (700, 12)); -- offset LSB 652
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s7173 => state := s7174;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (701, 12)); -- offset MSB 653
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7174 => state := s7175; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7175 => 			--4
	if (fixed2floatrdy = '1') then state := s7176;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7175; end if;
when s7176 => state := s7177; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7177 => 			--6
	if (mulfprdy = '1') then state := s7178;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7177; end if;
when s7178 => state := s7179; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7179 => 			--8
	if (mulfprdy = '1') then state := s7180;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7179; end if;
when s7180 => state := s7181; 	--9
	mulfpsclr <= '0';
when s7181 => state := s7182; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7182 => 			--11
	if (mulfprdy = '1') then state := s7183;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7182; end if;
when s7183 => state := s7184; 	--12
	mulfpsclr <= '0';
when s7184 => state := s7185; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7185 => 			--14
	if (addfprdy = '1') then state := s7186;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7185; end if;
when s7186 => state := s7187; 	--15
	addfpsclr <= '0';
when s7187 => state := s7188; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7188 => 			--17
	if (addfprdy = '1') then state := s7189;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7188; end if;
when s7189 => state := s7190; 	--18
	addfpsclr <= '0';
when s7190 => state := s7191; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7191 => 			--20
	if (addfprdy = '1') then state := s7192;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7191; end if;
when s7192 => state := s7193; 	--21
	addfpsclr <= '0';
when s7193 => state := s7194; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (382, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7194 => state := s7195; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (702, 12)); -- offset LSB 654
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s7195 => state := s7196;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (703, 12)); -- offset MSB 655
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7196 => state := s7197; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7197 => 			--4
	if (fixed2floatrdy = '1') then state := s7198;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7197; end if;
when s7198 => state := s7199; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7199 => 			--6
	if (mulfprdy = '1') then state := s7200;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7199; end if;
when s7200 => state := s7201; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7201 => 			--8
	if (mulfprdy = '1') then state := s7202;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7201; end if;
when s7202 => state := s7203; 	--9
	mulfpsclr <= '0';
when s7203 => state := s7204; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7204 => 			--11
	if (mulfprdy = '1') then state := s7205;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7204; end if;
when s7205 => state := s7206; 	--12
	mulfpsclr <= '0';
when s7206 => state := s7207; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7207 => 			--14
	if (addfprdy = '1') then state := s7208;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7207; end if;
when s7208 => state := s7209; 	--15
	addfpsclr <= '0';
when s7209 => state := s7210; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7210 => 			--17
	if (addfprdy = '1') then state := s7211;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7210; end if;
when s7211 => state := s7212; 	--18
	addfpsclr <= '0';
when s7212 => state := s7213; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7213 => 			--20
	if (addfprdy = '1') then state := s7214;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7213; end if;
when s7214 => state := s7215; 	--21
	addfpsclr <= '0';
when s7215 => state := s7216; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (383, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7216 => state := s7217; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (704, 12)); -- offset LSB 656
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s7217 => state := s7218;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (705, 12)); -- offset MSB 657
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7218 => state := s7219; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7219 => 			--4
	if (fixed2floatrdy = '1') then state := s7220;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7219; end if;
when s7220 => state := s7221; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7221 => 			--6
	if (mulfprdy = '1') then state := s7222;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7221; end if;
when s7222 => state := s7223; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7223 => 			--8
	if (mulfprdy = '1') then state := s7224;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7223; end if;
when s7224 => state := s7225; 	--9
	mulfpsclr <= '0';
when s7225 => state := s7226; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7226 => 			--11
	if (mulfprdy = '1') then state := s7227;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7226; end if;
when s7227 => state := s7228; 	--12
	mulfpsclr <= '0';
when s7228 => state := s7229; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7229 => 			--14
	if (addfprdy = '1') then state := s7230;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7229; end if;
when s7230 => state := s7231; 	--15
	addfpsclr <= '0';
when s7231 => state := s7232; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7232 => 			--17
	if (addfprdy = '1') then state := s7233;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7232; end if;
when s7233 => state := s7234; 	--18
	addfpsclr <= '0';
when s7234 => state := s7235; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7235 => 			--20
	if (addfprdy = '1') then state := s7236;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7235; end if;
when s7236 => state := s7237; 	--21
	addfpsclr <= '0';
when s7237 => state := s7238; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (384, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7238 => state := s7239; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (706, 12)); -- offset LSB 658
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s7239 => state := s7240;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (707, 12)); -- offset MSB 659
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7240 => state := s7241; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7241 => 			--4
	if (fixed2floatrdy = '1') then state := s7242;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7241; end if;
when s7242 => state := s7243; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7243 => 			--6
	if (mulfprdy = '1') then state := s7244;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7243; end if;
when s7244 => state := s7245; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7245 => 			--8
	if (mulfprdy = '1') then state := s7246;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7245; end if;
when s7246 => state := s7247; 	--9
	mulfpsclr <= '0';
when s7247 => state := s7248; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7248 => 			--11
	if (mulfprdy = '1') then state := s7249;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7248; end if;
when s7249 => state := s7250; 	--12
	mulfpsclr <= '0';
when s7250 => state := s7251; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7251 => 			--14
	if (addfprdy = '1') then state := s7252;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7251; end if;
when s7252 => state := s7253; 	--15
	addfpsclr <= '0';
when s7253 => state := s7254; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7254 => 			--17
	if (addfprdy = '1') then state := s7255;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7254; end if;
when s7255 => state := s7256; 	--18
	addfpsclr <= '0';
when s7256 => state := s7257; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7257 => 			--20
	if (addfprdy = '1') then state := s7258;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7257; end if;
when s7258 => state := s7259; 	--21
	addfpsclr <= '0';
when s7259 => state := s7260; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (385, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7260 => state := s7261; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (708, 12)); -- offset LSB 660
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s7261 => state := s7262;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (709, 12)); -- offset MSB 661
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7262 => state := s7263; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7263 => 			--4
	if (fixed2floatrdy = '1') then state := s7264;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7263; end if;
when s7264 => state := s7265; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7265 => 			--6
	if (mulfprdy = '1') then state := s7266;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7265; end if;
when s7266 => state := s7267; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7267 => 			--8
	if (mulfprdy = '1') then state := s7268;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7267; end if;
when s7268 => state := s7269; 	--9
	mulfpsclr <= '0';
when s7269 => state := s7270; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7270 => 			--11
	if (mulfprdy = '1') then state := s7271;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7270; end if;
when s7271 => state := s7272; 	--12
	mulfpsclr <= '0';
when s7272 => state := s7273; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7273 => 			--14
	if (addfprdy = '1') then state := s7274;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7273; end if;
when s7274 => state := s7275; 	--15
	addfpsclr <= '0';
when s7275 => state := s7276; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7276 => 			--17
	if (addfprdy = '1') then state := s7277;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7276; end if;
when s7277 => state := s7278; 	--18
	addfpsclr <= '0';
when s7278 => state := s7279; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7279 => 			--20
	if (addfprdy = '1') then state := s7280;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7279; end if;
when s7280 => state := s7281; 	--21
	addfpsclr <= '0';
when s7281 => state := s7282; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (386, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7282 => state := s7283; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (710, 12)); -- offset LSB 662
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s7283 => state := s7284;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (711, 12)); -- offset MSB 663
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7284 => state := s7285; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7285 => 			--4
	if (fixed2floatrdy = '1') then state := s7286;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7285; end if;
when s7286 => state := s7287; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7287 => 			--6
	if (mulfprdy = '1') then state := s7288;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7287; end if;
when s7288 => state := s7289; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7289 => 			--8
	if (mulfprdy = '1') then state := s7290;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7289; end if;
when s7290 => state := s7291; 	--9
	mulfpsclr <= '0';
when s7291 => state := s7292; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7292 => 			--11
	if (mulfprdy = '1') then state := s7293;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7292; end if;
when s7293 => state := s7294; 	--12
	mulfpsclr <= '0';
when s7294 => state := s7295; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7295 => 			--14
	if (addfprdy = '1') then state := s7296;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7295; end if;
when s7296 => state := s7297; 	--15
	addfpsclr <= '0';
when s7297 => state := s7298; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7298 => 			--17
	if (addfprdy = '1') then state := s7299;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7298; end if;
when s7299 => state := s7300; 	--18
	addfpsclr <= '0';
when s7300 => state := s7301; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7301 => 			--20
	if (addfprdy = '1') then state := s7302;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7301; end if;
when s7302 => state := s7303; 	--21
	addfpsclr <= '0';
when s7303 => state := s7304; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (387, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7304 => state := s7305; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (712, 12)); -- offset LSB 664
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s7305 => state := s7306;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (713, 12)); -- offset MSB 665
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7306 => state := s7307; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7307 => 			--4
	if (fixed2floatrdy = '1') then state := s7308;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7307; end if;
when s7308 => state := s7309; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7309 => 			--6
	if (mulfprdy = '1') then state := s7310;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7309; end if;
when s7310 => state := s7311; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7311 => 			--8
	if (mulfprdy = '1') then state := s7312;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7311; end if;
when s7312 => state := s7313; 	--9
	mulfpsclr <= '0';
when s7313 => state := s7314; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7314 => 			--11
	if (mulfprdy = '1') then state := s7315;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7314; end if;
when s7315 => state := s7316; 	--12
	mulfpsclr <= '0';
when s7316 => state := s7317; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7317 => 			--14
	if (addfprdy = '1') then state := s7318;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7317; end if;
when s7318 => state := s7319; 	--15
	addfpsclr <= '0';
when s7319 => state := s7320; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7320 => 			--17
	if (addfprdy = '1') then state := s7321;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7320; end if;
when s7321 => state := s7322; 	--18
	addfpsclr <= '0';
when s7322 => state := s7323; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7323 => 			--20
	if (addfprdy = '1') then state := s7324;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7323; end if;
when s7324 => state := s7325; 	--21
	addfpsclr <= '0';
when s7325 => state := s7326; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (388, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7326 => state := s7327; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (714, 12)); -- offset LSB 666
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s7327 => state := s7328;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (715, 12)); -- offset MSB 667
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7328 => state := s7329; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7329 => 			--4
	if (fixed2floatrdy = '1') then state := s7330;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7329; end if;
when s7330 => state := s7331; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7331 => 			--6
	if (mulfprdy = '1') then state := s7332;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7331; end if;
when s7332 => state := s7333; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7333 => 			--8
	if (mulfprdy = '1') then state := s7334;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7333; end if;
when s7334 => state := s7335; 	--9
	mulfpsclr <= '0';
when s7335 => state := s7336; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7336 => 			--11
	if (mulfprdy = '1') then state := s7337;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7336; end if;
when s7337 => state := s7338; 	--12
	mulfpsclr <= '0';
when s7338 => state := s7339; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7339 => 			--14
	if (addfprdy = '1') then state := s7340;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7339; end if;
when s7340 => state := s7341; 	--15
	addfpsclr <= '0';
when s7341 => state := s7342; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7342 => 			--17
	if (addfprdy = '1') then state := s7343;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7342; end if;
when s7343 => state := s7344; 	--18
	addfpsclr <= '0';
when s7344 => state := s7345; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7345 => 			--20
	if (addfprdy = '1') then state := s7346;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7345; end if;
when s7346 => state := s7347; 	--21
	addfpsclr <= '0';
when s7347 => state := s7348; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (389, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7348 => state := s7349; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (716, 12)); -- offset LSB 668
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s7349 => state := s7350;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (717, 12)); -- offset MSB 669
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7350 => state := s7351; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7351 => 			--4
	if (fixed2floatrdy = '1') then state := s7352;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7351; end if;
when s7352 => state := s7353; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7353 => 			--6
	if (mulfprdy = '1') then state := s7354;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7353; end if;
when s7354 => state := s7355; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7355 => 			--8
	if (mulfprdy = '1') then state := s7356;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7355; end if;
when s7356 => state := s7357; 	--9
	mulfpsclr <= '0';
when s7357 => state := s7358; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7358 => 			--11
	if (mulfprdy = '1') then state := s7359;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7358; end if;
when s7359 => state := s7360; 	--12
	mulfpsclr <= '0';
when s7360 => state := s7361; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7361 => 			--14
	if (addfprdy = '1') then state := s7362;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7361; end if;
when s7362 => state := s7363; 	--15
	addfpsclr <= '0';
when s7363 => state := s7364; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7364 => 			--17
	if (addfprdy = '1') then state := s7365;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7364; end if;
when s7365 => state := s7366; 	--18
	addfpsclr <= '0';
when s7366 => state := s7367; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7367 => 			--20
	if (addfprdy = '1') then state := s7368;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7367; end if;
when s7368 => state := s7369; 	--21
	addfpsclr <= '0';
when s7369 => state := s7370; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (390, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7370 => state := s7371; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (718, 12)); -- offset LSB 670
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s7371 => state := s7372;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (719, 12)); -- offset MSB 671
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7372 => state := s7373; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7373 => 			--4
	if (fixed2floatrdy = '1') then state := s7374;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7373; end if;
when s7374 => state := s7375; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7375 => 			--6
	if (mulfprdy = '1') then state := s7376;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7375; end if;
when s7376 => state := s7377; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7377 => 			--8
	if (mulfprdy = '1') then state := s7378;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7377; end if;
when s7378 => state := s7379; 	--9
	mulfpsclr <= '0';
when s7379 => state := s7380; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7380 => 			--11
	if (mulfprdy = '1') then state := s7381;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7380; end if;
when s7381 => state := s7382; 	--12
	mulfpsclr <= '0';
when s7382 => state := s7383; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7383 => 			--14
	if (addfprdy = '1') then state := s7384;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7383; end if;
when s7384 => state := s7385; 	--15
	addfpsclr <= '0';
when s7385 => state := s7386; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7386 => 			--17
	if (addfprdy = '1') then state := s7387;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7386; end if;
when s7387 => state := s7388; 	--18
	addfpsclr <= '0';
when s7388 => state := s7389; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7389 => 			--20
	if (addfprdy = '1') then state := s7390;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7389; end if;
when s7390 => state := s7391; 	--21
	addfpsclr <= '0';
when s7391 => state := s7392; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (391, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7392 => state := s7393; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (720, 12)); -- offset LSB 672
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s7393 => state := s7394;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (721, 12)); -- offset MSB 673
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7394 => state := s7395; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7395 => 			--4
	if (fixed2floatrdy = '1') then state := s7396;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7395; end if;
when s7396 => state := s7397; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7397 => 			--6
	if (mulfprdy = '1') then state := s7398;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7397; end if;
when s7398 => state := s7399; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7399 => 			--8
	if (mulfprdy = '1') then state := s7400;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7399; end if;
when s7400 => state := s7401; 	--9
	mulfpsclr <= '0';
when s7401 => state := s7402; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7402 => 			--11
	if (mulfprdy = '1') then state := s7403;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7402; end if;
when s7403 => state := s7404; 	--12
	mulfpsclr <= '0';
when s7404 => state := s7405; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7405 => 			--14
	if (addfprdy = '1') then state := s7406;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7405; end if;
when s7406 => state := s7407; 	--15
	addfpsclr <= '0';
when s7407 => state := s7408; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7408 => 			--17
	if (addfprdy = '1') then state := s7409;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7408; end if;
when s7409 => state := s7410; 	--18
	addfpsclr <= '0';
when s7410 => state := s7411; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7411 => 			--20
	if (addfprdy = '1') then state := s7412;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7411; end if;
when s7412 => state := s7413; 	--21
	addfpsclr <= '0';
when s7413 => state := s7414; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (392, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7414 => state := s7415; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (722, 12)); -- offset LSB 674
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s7415 => state := s7416;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (723, 12)); -- offset MSB 675
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7416 => state := s7417; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7417 => 			--4
	if (fixed2floatrdy = '1') then state := s7418;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7417; end if;
when s7418 => state := s7419; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7419 => 			--6
	if (mulfprdy = '1') then state := s7420;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7419; end if;
when s7420 => state := s7421; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7421 => 			--8
	if (mulfprdy = '1') then state := s7422;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7421; end if;
when s7422 => state := s7423; 	--9
	mulfpsclr <= '0';
when s7423 => state := s7424; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7424 => 			--11
	if (mulfprdy = '1') then state := s7425;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7424; end if;
when s7425 => state := s7426; 	--12
	mulfpsclr <= '0';
when s7426 => state := s7427; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7427 => 			--14
	if (addfprdy = '1') then state := s7428;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7427; end if;
when s7428 => state := s7429; 	--15
	addfpsclr <= '0';
when s7429 => state := s7430; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7430 => 			--17
	if (addfprdy = '1') then state := s7431;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7430; end if;
when s7431 => state := s7432; 	--18
	addfpsclr <= '0';
when s7432 => state := s7433; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7433 => 			--20
	if (addfprdy = '1') then state := s7434;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7433; end if;
when s7434 => state := s7435; 	--21
	addfpsclr <= '0';
when s7435 => state := s7436; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (393, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7436 => state := s7437; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (724, 12)); -- offset LSB 676
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s7437 => state := s7438;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (725, 12)); -- offset MSB 677
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7438 => state := s7439; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7439 => 			--4
	if (fixed2floatrdy = '1') then state := s7440;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7439; end if;
when s7440 => state := s7441; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7441 => 			--6
	if (mulfprdy = '1') then state := s7442;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7441; end if;
when s7442 => state := s7443; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7443 => 			--8
	if (mulfprdy = '1') then state := s7444;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7443; end if;
when s7444 => state := s7445; 	--9
	mulfpsclr <= '0';
when s7445 => state := s7446; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7446 => 			--11
	if (mulfprdy = '1') then state := s7447;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7446; end if;
when s7447 => state := s7448; 	--12
	mulfpsclr <= '0';
when s7448 => state := s7449; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7449 => 			--14
	if (addfprdy = '1') then state := s7450;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7449; end if;
when s7450 => state := s7451; 	--15
	addfpsclr <= '0';
when s7451 => state := s7452; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7452 => 			--17
	if (addfprdy = '1') then state := s7453;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7452; end if;
when s7453 => state := s7454; 	--18
	addfpsclr <= '0';
when s7454 => state := s7455; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7455 => 			--20
	if (addfprdy = '1') then state := s7456;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7455; end if;
when s7456 => state := s7457; 	--21
	addfpsclr <= '0';
when s7457 => state := s7458; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (394, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7458 => state := s7459; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (726, 12)); -- offset LSB 678
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s7459 => state := s7460;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (727, 12)); -- offset MSB 679
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7460 => state := s7461; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7461 => 			--4
	if (fixed2floatrdy = '1') then state := s7462;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7461; end if;
when s7462 => state := s7463; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7463 => 			--6
	if (mulfprdy = '1') then state := s7464;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7463; end if;
when s7464 => state := s7465; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7465 => 			--8
	if (mulfprdy = '1') then state := s7466;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7465; end if;
when s7466 => state := s7467; 	--9
	mulfpsclr <= '0';
when s7467 => state := s7468; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7468 => 			--11
	if (mulfprdy = '1') then state := s7469;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7468; end if;
when s7469 => state := s7470; 	--12
	mulfpsclr <= '0';
when s7470 => state := s7471; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7471 => 			--14
	if (addfprdy = '1') then state := s7472;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7471; end if;
when s7472 => state := s7473; 	--15
	addfpsclr <= '0';
when s7473 => state := s7474; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7474 => 			--17
	if (addfprdy = '1') then state := s7475;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7474; end if;
when s7475 => state := s7476; 	--18
	addfpsclr <= '0';
when s7476 => state := s7477; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7477 => 			--20
	if (addfprdy = '1') then state := s7478;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7477; end if;
when s7478 => state := s7479; 	--21
	addfpsclr <= '0';
when s7479 => state := s7480; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (395, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7480 => state := s7481; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (728, 12)); -- offset LSB 680
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s7481 => state := s7482;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (729, 12)); -- offset MSB 681
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7482 => state := s7483; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7483 => 			--4
	if (fixed2floatrdy = '1') then state := s7484;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7483; end if;
when s7484 => state := s7485; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7485 => 			--6
	if (mulfprdy = '1') then state := s7486;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7485; end if;
when s7486 => state := s7487; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7487 => 			--8
	if (mulfprdy = '1') then state := s7488;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7487; end if;
when s7488 => state := s7489; 	--9
	mulfpsclr <= '0';
when s7489 => state := s7490; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7490 => 			--11
	if (mulfprdy = '1') then state := s7491;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7490; end if;
when s7491 => state := s7492; 	--12
	mulfpsclr <= '0';
when s7492 => state := s7493; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7493 => 			--14
	if (addfprdy = '1') then state := s7494;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7493; end if;
when s7494 => state := s7495; 	--15
	addfpsclr <= '0';
when s7495 => state := s7496; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7496 => 			--17
	if (addfprdy = '1') then state := s7497;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7496; end if;
when s7497 => state := s7498; 	--18
	addfpsclr <= '0';
when s7498 => state := s7499; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7499 => 			--20
	if (addfprdy = '1') then state := s7500;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7499; end if;
when s7500 => state := s7501; 	--21
	addfpsclr <= '0';
when s7501 => state := s7502; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (396, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7502 => state := s7503; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (730, 12)); -- offset LSB 682
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s7503 => state := s7504;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (731, 12)); -- offset MSB 683
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7504 => state := s7505; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7505 => 			--4
	if (fixed2floatrdy = '1') then state := s7506;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7505; end if;
when s7506 => state := s7507; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7507 => 			--6
	if (mulfprdy = '1') then state := s7508;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7507; end if;
when s7508 => state := s7509; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7509 => 			--8
	if (mulfprdy = '1') then state := s7510;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7509; end if;
when s7510 => state := s7511; 	--9
	mulfpsclr <= '0';
when s7511 => state := s7512; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7512 => 			--11
	if (mulfprdy = '1') then state := s7513;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7512; end if;
when s7513 => state := s7514; 	--12
	mulfpsclr <= '0';
when s7514 => state := s7515; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7515 => 			--14
	if (addfprdy = '1') then state := s7516;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7515; end if;
when s7516 => state := s7517; 	--15
	addfpsclr <= '0';
when s7517 => state := s7518; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7518 => 			--17
	if (addfprdy = '1') then state := s7519;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7518; end if;
when s7519 => state := s7520; 	--18
	addfpsclr <= '0';
when s7520 => state := s7521; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7521 => 			--20
	if (addfprdy = '1') then state := s7522;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7521; end if;
when s7522 => state := s7523; 	--21
	addfpsclr <= '0';
when s7523 => state := s7524; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (397, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7524 => state := s7525; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (732, 12)); -- offset LSB 684
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s7525 => state := s7526;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (733, 12)); -- offset MSB 685
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7526 => state := s7527; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7527 => 			--4
	if (fixed2floatrdy = '1') then state := s7528;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7527; end if;
when s7528 => state := s7529; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7529 => 			--6
	if (mulfprdy = '1') then state := s7530;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7529; end if;
when s7530 => state := s7531; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7531 => 			--8
	if (mulfprdy = '1') then state := s7532;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7531; end if;
when s7532 => state := s7533; 	--9
	mulfpsclr <= '0';
when s7533 => state := s7534; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7534 => 			--11
	if (mulfprdy = '1') then state := s7535;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7534; end if;
when s7535 => state := s7536; 	--12
	mulfpsclr <= '0';
when s7536 => state := s7537; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7537 => 			--14
	if (addfprdy = '1') then state := s7538;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7537; end if;
when s7538 => state := s7539; 	--15
	addfpsclr <= '0';
when s7539 => state := s7540; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7540 => 			--17
	if (addfprdy = '1') then state := s7541;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7540; end if;
when s7541 => state := s7542; 	--18
	addfpsclr <= '0';
when s7542 => state := s7543; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7543 => 			--20
	if (addfprdy = '1') then state := s7544;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7543; end if;
when s7544 => state := s7545; 	--21
	addfpsclr <= '0';
when s7545 => state := s7546; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (398, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7546 => state := s7547; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (734, 12)); -- offset LSB 686
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s7547 => state := s7548;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (735, 12)); -- offset MSB 687
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7548 => state := s7549; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7549 => 			--4
	if (fixed2floatrdy = '1') then state := s7550;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7549; end if;
when s7550 => state := s7551; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7551 => 			--6
	if (mulfprdy = '1') then state := s7552;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7551; end if;
when s7552 => state := s7553; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7553 => 			--8
	if (mulfprdy = '1') then state := s7554;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7553; end if;
when s7554 => state := s7555; 	--9
	mulfpsclr <= '0';
when s7555 => state := s7556; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7556 => 			--11
	if (mulfprdy = '1') then state := s7557;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7556; end if;
when s7557 => state := s7558; 	--12
	mulfpsclr <= '0';
when s7558 => state := s7559; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7559 => 			--14
	if (addfprdy = '1') then state := s7560;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7559; end if;
when s7560 => state := s7561; 	--15
	addfpsclr <= '0';
when s7561 => state := s7562; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7562 => 			--17
	if (addfprdy = '1') then state := s7563;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7562; end if;
when s7563 => state := s7564; 	--18
	addfpsclr <= '0';
when s7564 => state := s7565; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7565 => 			--20
	if (addfprdy = '1') then state := s7566;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7565; end if;
when s7566 => state := s7567; 	--21
	addfpsclr <= '0';
when s7567 => state := s7568; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (399, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7568 => state := s7569; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (736, 12)); -- offset LSB 688
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s7569 => state := s7570;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (737, 12)); -- offset MSB 689
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7570 => state := s7571; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7571 => 			--4
	if (fixed2floatrdy = '1') then state := s7572;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7571; end if;
when s7572 => state := s7573; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7573 => 			--6
	if (mulfprdy = '1') then state := s7574;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7573; end if;
when s7574 => state := s7575; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7575 => 			--8
	if (mulfprdy = '1') then state := s7576;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7575; end if;
when s7576 => state := s7577; 	--9
	mulfpsclr <= '0';
when s7577 => state := s7578; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7578 => 			--11
	if (mulfprdy = '1') then state := s7579;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7578; end if;
when s7579 => state := s7580; 	--12
	mulfpsclr <= '0';
when s7580 => state := s7581; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7581 => 			--14
	if (addfprdy = '1') then state := s7582;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7581; end if;
when s7582 => state := s7583; 	--15
	addfpsclr <= '0';
when s7583 => state := s7584; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7584 => 			--17
	if (addfprdy = '1') then state := s7585;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7584; end if;
when s7585 => state := s7586; 	--18
	addfpsclr <= '0';
when s7586 => state := s7587; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7587 => 			--20
	if (addfprdy = '1') then state := s7588;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7587; end if;
when s7588 => state := s7589; 	--21
	addfpsclr <= '0';
when s7589 => state := s7590; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (400, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7590 => state := s7591; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (738, 12)); -- offset LSB 690
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s7591 => state := s7592;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (739, 12)); -- offset MSB 691
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7592 => state := s7593; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7593 => 			--4
	if (fixed2floatrdy = '1') then state := s7594;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7593; end if;
when s7594 => state := s7595; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7595 => 			--6
	if (mulfprdy = '1') then state := s7596;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7595; end if;
when s7596 => state := s7597; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7597 => 			--8
	if (mulfprdy = '1') then state := s7598;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7597; end if;
when s7598 => state := s7599; 	--9
	mulfpsclr <= '0';
when s7599 => state := s7600; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7600 => 			--11
	if (mulfprdy = '1') then state := s7601;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7600; end if;
when s7601 => state := s7602; 	--12
	mulfpsclr <= '0';
when s7602 => state := s7603; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7603 => 			--14
	if (addfprdy = '1') then state := s7604;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7603; end if;
when s7604 => state := s7605; 	--15
	addfpsclr <= '0';
when s7605 => state := s7606; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7606 => 			--17
	if (addfprdy = '1') then state := s7607;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7606; end if;
when s7607 => state := s7608; 	--18
	addfpsclr <= '0';
when s7608 => state := s7609; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7609 => 			--20
	if (addfprdy = '1') then state := s7610;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7609; end if;
when s7610 => state := s7611; 	--21
	addfpsclr <= '0';
when s7611 => state := s7612; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (401, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7612 => state := s7613; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (740, 12)); -- offset LSB 692
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s7613 => state := s7614;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (741, 12)); -- offset MSB 693
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7614 => state := s7615; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7615 => 			--4
	if (fixed2floatrdy = '1') then state := s7616;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7615; end if;
when s7616 => state := s7617; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7617 => 			--6
	if (mulfprdy = '1') then state := s7618;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7617; end if;
when s7618 => state := s7619; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7619 => 			--8
	if (mulfprdy = '1') then state := s7620;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7619; end if;
when s7620 => state := s7621; 	--9
	mulfpsclr <= '0';
when s7621 => state := s7622; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7622 => 			--11
	if (mulfprdy = '1') then state := s7623;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7622; end if;
when s7623 => state := s7624; 	--12
	mulfpsclr <= '0';
when s7624 => state := s7625; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7625 => 			--14
	if (addfprdy = '1') then state := s7626;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7625; end if;
when s7626 => state := s7627; 	--15
	addfpsclr <= '0';
when s7627 => state := s7628; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7628 => 			--17
	if (addfprdy = '1') then state := s7629;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7628; end if;
when s7629 => state := s7630; 	--18
	addfpsclr <= '0';
when s7630 => state := s7631; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7631 => 			--20
	if (addfprdy = '1') then state := s7632;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7631; end if;
when s7632 => state := s7633; 	--21
	addfpsclr <= '0';
when s7633 => state := s7634; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (402, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7634 => state := s7635; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (742, 12)); -- offset LSB 694
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s7635 => state := s7636;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (743, 12)); -- offset MSB 695
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7636 => state := s7637; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7637 => 			--4
	if (fixed2floatrdy = '1') then state := s7638;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7637; end if;
when s7638 => state := s7639; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7639 => 			--6
	if (mulfprdy = '1') then state := s7640;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7639; end if;
when s7640 => state := s7641; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7641 => 			--8
	if (mulfprdy = '1') then state := s7642;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7641; end if;
when s7642 => state := s7643; 	--9
	mulfpsclr <= '0';
when s7643 => state := s7644; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7644 => 			--11
	if (mulfprdy = '1') then state := s7645;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7644; end if;
when s7645 => state := s7646; 	--12
	mulfpsclr <= '0';
when s7646 => state := s7647; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7647 => 			--14
	if (addfprdy = '1') then state := s7648;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7647; end if;
when s7648 => state := s7649; 	--15
	addfpsclr <= '0';
when s7649 => state := s7650; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7650 => 			--17
	if (addfprdy = '1') then state := s7651;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7650; end if;
when s7651 => state := s7652; 	--18
	addfpsclr <= '0';
when s7652 => state := s7653; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7653 => 			--20
	if (addfprdy = '1') then state := s7654;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7653; end if;
when s7654 => state := s7655; 	--21
	addfpsclr <= '0';
when s7655 => state := s7656; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (403, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7656 => state := s7657; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (744, 12)); -- offset LSB 696
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s7657 => state := s7658;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (745, 12)); -- offset MSB 697
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7658 => state := s7659; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7659 => 			--4
	if (fixed2floatrdy = '1') then state := s7660;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7659; end if;
when s7660 => state := s7661; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7661 => 			--6
	if (mulfprdy = '1') then state := s7662;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7661; end if;
when s7662 => state := s7663; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7663 => 			--8
	if (mulfprdy = '1') then state := s7664;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7663; end if;
when s7664 => state := s7665; 	--9
	mulfpsclr <= '0';
when s7665 => state := s7666; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7666 => 			--11
	if (mulfprdy = '1') then state := s7667;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7666; end if;
when s7667 => state := s7668; 	--12
	mulfpsclr <= '0';
when s7668 => state := s7669; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7669 => 			--14
	if (addfprdy = '1') then state := s7670;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7669; end if;
when s7670 => state := s7671; 	--15
	addfpsclr <= '0';
when s7671 => state := s7672; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7672 => 			--17
	if (addfprdy = '1') then state := s7673;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7672; end if;
when s7673 => state := s7674; 	--18
	addfpsclr <= '0';
when s7674 => state := s7675; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7675 => 			--20
	if (addfprdy = '1') then state := s7676;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7675; end if;
when s7676 => state := s7677; 	--21
	addfpsclr <= '0';
when s7677 => state := s7678; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (404, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7678 => state := s7679; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (746, 12)); -- offset LSB 698
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s7679 => state := s7680;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (747, 12)); -- offset MSB 699
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7680 => state := s7681; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7681 => 			--4
	if (fixed2floatrdy = '1') then state := s7682;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7681; end if;
when s7682 => state := s7683; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7683 => 			--6
	if (mulfprdy = '1') then state := s7684;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7683; end if;
when s7684 => state := s7685; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7685 => 			--8
	if (mulfprdy = '1') then state := s7686;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7685; end if;
when s7686 => state := s7687; 	--9
	mulfpsclr <= '0';
when s7687 => state := s7688; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7688 => 			--11
	if (mulfprdy = '1') then state := s7689;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7688; end if;
when s7689 => state := s7690; 	--12
	mulfpsclr <= '0';
when s7690 => state := s7691; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7691 => 			--14
	if (addfprdy = '1') then state := s7692;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7691; end if;
when s7692 => state := s7693; 	--15
	addfpsclr <= '0';
when s7693 => state := s7694; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7694 => 			--17
	if (addfprdy = '1') then state := s7695;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7694; end if;
when s7695 => state := s7696; 	--18
	addfpsclr <= '0';
when s7696 => state := s7697; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7697 => 			--20
	if (addfprdy = '1') then state := s7698;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7697; end if;
when s7698 => state := s7699; 	--21
	addfpsclr <= '0';
when s7699 => state := s7700; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (405, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7700 => state := s7701; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (748, 12)); -- offset LSB 700
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s7701 => state := s7702;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (749, 12)); -- offset MSB 701
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7702 => state := s7703; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7703 => 			--4
	if (fixed2floatrdy = '1') then state := s7704;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7703; end if;
when s7704 => state := s7705; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7705 => 			--6
	if (mulfprdy = '1') then state := s7706;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7705; end if;
when s7706 => state := s7707; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7707 => 			--8
	if (mulfprdy = '1') then state := s7708;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7707; end if;
when s7708 => state := s7709; 	--9
	mulfpsclr <= '0';
when s7709 => state := s7710; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7710 => 			--11
	if (mulfprdy = '1') then state := s7711;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7710; end if;
when s7711 => state := s7712; 	--12
	mulfpsclr <= '0';
when s7712 => state := s7713; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7713 => 			--14
	if (addfprdy = '1') then state := s7714;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7713; end if;
when s7714 => state := s7715; 	--15
	addfpsclr <= '0';
when s7715 => state := s7716; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7716 => 			--17
	if (addfprdy = '1') then state := s7717;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7716; end if;
when s7717 => state := s7718; 	--18
	addfpsclr <= '0';
when s7718 => state := s7719; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7719 => 			--20
	if (addfprdy = '1') then state := s7720;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7719; end if;
when s7720 => state := s7721; 	--21
	addfpsclr <= '0';
when s7721 => state := s7722; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (406, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7722 => state := s7723; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (750, 12)); -- offset LSB 702
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s7723 => state := s7724;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (751, 12)); -- offset MSB 703
	addra <= std_logic_vector (to_unsigned (10, 10)); -- OCCrowI 10
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7724 => state := s7725; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7725 => 			--4
	if (fixed2floatrdy = '1') then state := s7726;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7725; end if;
when s7726 => state := s7727; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7727 => 			--6
	if (mulfprdy = '1') then state := s7728;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7727; end if;
when s7728 => state := s7729; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7729 => 			--8
	if (mulfprdy = '1') then state := s7730;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7729; end if;
when s7730 => state := s7731; 	--9
	mulfpsclr <= '0';
when s7731 => state := s7732; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7732 => 			--11
	if (mulfprdy = '1') then state := s7733;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7732; end if;
when s7733 => state := s7734; 	--12
	mulfpsclr <= '0';
when s7734 => state := s7735; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7735 => 			--14
	if (addfprdy = '1') then state := s7736;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7735; end if;
when s7736 => state := s7737; 	--15
	addfpsclr <= '0';
when s7737 => state := s7738; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7738 => 			--17
	if (addfprdy = '1') then state := s7739;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7738; end if;
when s7739 => state := s7740; 	--18
	addfpsclr <= '0';
when s7740 => state := s7741; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7741 => 			--20
	if (addfprdy = '1') then state := s7742;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7741; end if;
when s7742 => state := s7743; 	--21
	addfpsclr <= '0';
when s7743 => state := s7744; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (407, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7744 => state := s7745; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (752, 12)); -- offset LSB 704
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s7745 => state := s7746;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (753, 12)); -- offset MSB 705
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7746 => state := s7747; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7747 => 			--4
	if (fixed2floatrdy = '1') then state := s7748;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7747; end if;
when s7748 => state := s7749; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7749 => 			--6
	if (mulfprdy = '1') then state := s7750;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7749; end if;
when s7750 => state := s7751; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7751 => 			--8
	if (mulfprdy = '1') then state := s7752;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7751; end if;
when s7752 => state := s7753; 	--9
	mulfpsclr <= '0';
when s7753 => state := s7754; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7754 => 			--11
	if (mulfprdy = '1') then state := s7755;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7754; end if;
when s7755 => state := s7756; 	--12
	mulfpsclr <= '0';
when s7756 => state := s7757; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7757 => 			--14
	if (addfprdy = '1') then state := s7758;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7757; end if;
when s7758 => state := s7759; 	--15
	addfpsclr <= '0';
when s7759 => state := s7760; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7760 => 			--17
	if (addfprdy = '1') then state := s7761;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7760; end if;
when s7761 => state := s7762; 	--18
	addfpsclr <= '0';
when s7762 => state := s7763; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7763 => 			--20
	if (addfprdy = '1') then state := s7764;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7763; end if;
when s7764 => state := s7765; 	--21
	addfpsclr <= '0';
when s7765 => state := s7766; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (408, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7766 => state := s7767; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (754, 12)); -- offset LSB 706
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s7767 => state := s7768;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (755, 12)); -- offset MSB 707
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7768 => state := s7769; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7769 => 			--4
	if (fixed2floatrdy = '1') then state := s7770;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7769; end if;
when s7770 => state := s7771; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7771 => 			--6
	if (mulfprdy = '1') then state := s7772;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7771; end if;
when s7772 => state := s7773; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7773 => 			--8
	if (mulfprdy = '1') then state := s7774;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7773; end if;
when s7774 => state := s7775; 	--9
	mulfpsclr <= '0';
when s7775 => state := s7776; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7776 => 			--11
	if (mulfprdy = '1') then state := s7777;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7776; end if;
when s7777 => state := s7778; 	--12
	mulfpsclr <= '0';
when s7778 => state := s7779; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7779 => 			--14
	if (addfprdy = '1') then state := s7780;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7779; end if;
when s7780 => state := s7781; 	--15
	addfpsclr <= '0';
when s7781 => state := s7782; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7782 => 			--17
	if (addfprdy = '1') then state := s7783;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7782; end if;
when s7783 => state := s7784; 	--18
	addfpsclr <= '0';
when s7784 => state := s7785; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7785 => 			--20
	if (addfprdy = '1') then state := s7786;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7785; end if;
when s7786 => state := s7787; 	--21
	addfpsclr <= '0';
when s7787 => state := s7788; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (409, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7788 => state := s7789; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (756, 12)); -- offset LSB 708
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s7789 => state := s7790;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (757, 12)); -- offset MSB 709
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7790 => state := s7791; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7791 => 			--4
	if (fixed2floatrdy = '1') then state := s7792;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7791; end if;
when s7792 => state := s7793; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7793 => 			--6
	if (mulfprdy = '1') then state := s7794;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7793; end if;
when s7794 => state := s7795; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7795 => 			--8
	if (mulfprdy = '1') then state := s7796;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7795; end if;
when s7796 => state := s7797; 	--9
	mulfpsclr <= '0';
when s7797 => state := s7798; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7798 => 			--11
	if (mulfprdy = '1') then state := s7799;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7798; end if;
when s7799 => state := s7800; 	--12
	mulfpsclr <= '0';
when s7800 => state := s7801; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7801 => 			--14
	if (addfprdy = '1') then state := s7802;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7801; end if;
when s7802 => state := s7803; 	--15
	addfpsclr <= '0';
when s7803 => state := s7804; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7804 => 			--17
	if (addfprdy = '1') then state := s7805;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7804; end if;
when s7805 => state := s7806; 	--18
	addfpsclr <= '0';
when s7806 => state := s7807; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7807 => 			--20
	if (addfprdy = '1') then state := s7808;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7807; end if;
when s7808 => state := s7809; 	--21
	addfpsclr <= '0';
when s7809 => state := s7810; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (410, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7810 => state := s7811; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (758, 12)); -- offset LSB 710
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s7811 => state := s7812;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (759, 12)); -- offset MSB 711
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7812 => state := s7813; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7813 => 			--4
	if (fixed2floatrdy = '1') then state := s7814;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7813; end if;
when s7814 => state := s7815; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7815 => 			--6
	if (mulfprdy = '1') then state := s7816;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7815; end if;
when s7816 => state := s7817; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7817 => 			--8
	if (mulfprdy = '1') then state := s7818;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7817; end if;
when s7818 => state := s7819; 	--9
	mulfpsclr <= '0';
when s7819 => state := s7820; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7820 => 			--11
	if (mulfprdy = '1') then state := s7821;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7820; end if;
when s7821 => state := s7822; 	--12
	mulfpsclr <= '0';
when s7822 => state := s7823; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7823 => 			--14
	if (addfprdy = '1') then state := s7824;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7823; end if;
when s7824 => state := s7825; 	--15
	addfpsclr <= '0';
when s7825 => state := s7826; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7826 => 			--17
	if (addfprdy = '1') then state := s7827;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7826; end if;
when s7827 => state := s7828; 	--18
	addfpsclr <= '0';
when s7828 => state := s7829; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7829 => 			--20
	if (addfprdy = '1') then state := s7830;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7829; end if;
when s7830 => state := s7831; 	--21
	addfpsclr <= '0';
when s7831 => state := s7832; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (411, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7832 => state := s7833; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (760, 12)); -- offset LSB 712
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s7833 => state := s7834;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (761, 12)); -- offset MSB 713
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7834 => state := s7835; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7835 => 			--4
	if (fixed2floatrdy = '1') then state := s7836;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7835; end if;
when s7836 => state := s7837; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7837 => 			--6
	if (mulfprdy = '1') then state := s7838;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7837; end if;
when s7838 => state := s7839; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7839 => 			--8
	if (mulfprdy = '1') then state := s7840;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7839; end if;
when s7840 => state := s7841; 	--9
	mulfpsclr <= '0';
when s7841 => state := s7842; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7842 => 			--11
	if (mulfprdy = '1') then state := s7843;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7842; end if;
when s7843 => state := s7844; 	--12
	mulfpsclr <= '0';
when s7844 => state := s7845; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7845 => 			--14
	if (addfprdy = '1') then state := s7846;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7845; end if;
when s7846 => state := s7847; 	--15
	addfpsclr <= '0';
when s7847 => state := s7848; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7848 => 			--17
	if (addfprdy = '1') then state := s7849;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7848; end if;
when s7849 => state := s7850; 	--18
	addfpsclr <= '0';
when s7850 => state := s7851; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7851 => 			--20
	if (addfprdy = '1') then state := s7852;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7851; end if;
when s7852 => state := s7853; 	--21
	addfpsclr <= '0';
when s7853 => state := s7854; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (412, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7854 => state := s7855; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (762, 12)); -- offset LSB 714
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s7855 => state := s7856;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (763, 12)); -- offset MSB 715
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7856 => state := s7857; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7857 => 			--4
	if (fixed2floatrdy = '1') then state := s7858;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7857; end if;
when s7858 => state := s7859; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7859 => 			--6
	if (mulfprdy = '1') then state := s7860;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7859; end if;
when s7860 => state := s7861; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7861 => 			--8
	if (mulfprdy = '1') then state := s7862;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7861; end if;
when s7862 => state := s7863; 	--9
	mulfpsclr <= '0';
when s7863 => state := s7864; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7864 => 			--11
	if (mulfprdy = '1') then state := s7865;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7864; end if;
when s7865 => state := s7866; 	--12
	mulfpsclr <= '0';
when s7866 => state := s7867; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7867 => 			--14
	if (addfprdy = '1') then state := s7868;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7867; end if;
when s7868 => state := s7869; 	--15
	addfpsclr <= '0';
when s7869 => state := s7870; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7870 => 			--17
	if (addfprdy = '1') then state := s7871;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7870; end if;
when s7871 => state := s7872; 	--18
	addfpsclr <= '0';
when s7872 => state := s7873; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7873 => 			--20
	if (addfprdy = '1') then state := s7874;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7873; end if;
when s7874 => state := s7875; 	--21
	addfpsclr <= '0';
when s7875 => state := s7876; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (413, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7876 => state := s7877; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (764, 12)); -- offset LSB 716
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s7877 => state := s7878;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (765, 12)); -- offset MSB 717
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7878 => state := s7879; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7879 => 			--4
	if (fixed2floatrdy = '1') then state := s7880;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7879; end if;
when s7880 => state := s7881; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7881 => 			--6
	if (mulfprdy = '1') then state := s7882;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7881; end if;
when s7882 => state := s7883; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7883 => 			--8
	if (mulfprdy = '1') then state := s7884;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7883; end if;
when s7884 => state := s7885; 	--9
	mulfpsclr <= '0';
when s7885 => state := s7886; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7886 => 			--11
	if (mulfprdy = '1') then state := s7887;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7886; end if;
when s7887 => state := s7888; 	--12
	mulfpsclr <= '0';
when s7888 => state := s7889; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7889 => 			--14
	if (addfprdy = '1') then state := s7890;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7889; end if;
when s7890 => state := s7891; 	--15
	addfpsclr <= '0';
when s7891 => state := s7892; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7892 => 			--17
	if (addfprdy = '1') then state := s7893;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7892; end if;
when s7893 => state := s7894; 	--18
	addfpsclr <= '0';
when s7894 => state := s7895; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7895 => 			--20
	if (addfprdy = '1') then state := s7896;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7895; end if;
when s7896 => state := s7897; 	--21
	addfpsclr <= '0';
when s7897 => state := s7898; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (414, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7898 => state := s7899; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (766, 12)); -- offset LSB 718
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s7899 => state := s7900;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (767, 12)); -- offset MSB 719
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7900 => state := s7901; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7901 => 			--4
	if (fixed2floatrdy = '1') then state := s7902;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7901; end if;
when s7902 => state := s7903; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7903 => 			--6
	if (mulfprdy = '1') then state := s7904;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7903; end if;
when s7904 => state := s7905; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7905 => 			--8
	if (mulfprdy = '1') then state := s7906;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7905; end if;
when s7906 => state := s7907; 	--9
	mulfpsclr <= '0';
when s7907 => state := s7908; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7908 => 			--11
	if (mulfprdy = '1') then state := s7909;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7908; end if;
when s7909 => state := s7910; 	--12
	mulfpsclr <= '0';
when s7910 => state := s7911; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7911 => 			--14
	if (addfprdy = '1') then state := s7912;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7911; end if;
when s7912 => state := s7913; 	--15
	addfpsclr <= '0';
when s7913 => state := s7914; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7914 => 			--17
	if (addfprdy = '1') then state := s7915;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7914; end if;
when s7915 => state := s7916; 	--18
	addfpsclr <= '0';
when s7916 => state := s7917; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7917 => 			--20
	if (addfprdy = '1') then state := s7918;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7917; end if;
when s7918 => state := s7919; 	--21
	addfpsclr <= '0';
when s7919 => state := s7920; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (415, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7920 => state := s7921; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (768, 12)); -- offset LSB 720
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s7921 => state := s7922;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (769, 12)); -- offset MSB 721
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7922 => state := s7923; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7923 => 			--4
	if (fixed2floatrdy = '1') then state := s7924;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7923; end if;
when s7924 => state := s7925; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7925 => 			--6
	if (mulfprdy = '1') then state := s7926;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7925; end if;
when s7926 => state := s7927; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7927 => 			--8
	if (mulfprdy = '1') then state := s7928;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7927; end if;
when s7928 => state := s7929; 	--9
	mulfpsclr <= '0';
when s7929 => state := s7930; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7930 => 			--11
	if (mulfprdy = '1') then state := s7931;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7930; end if;
when s7931 => state := s7932; 	--12
	mulfpsclr <= '0';
when s7932 => state := s7933; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7933 => 			--14
	if (addfprdy = '1') then state := s7934;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7933; end if;
when s7934 => state := s7935; 	--15
	addfpsclr <= '0';
when s7935 => state := s7936; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7936 => 			--17
	if (addfprdy = '1') then state := s7937;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7936; end if;
when s7937 => state := s7938; 	--18
	addfpsclr <= '0';
when s7938 => state := s7939; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7939 => 			--20
	if (addfprdy = '1') then state := s7940;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7939; end if;
when s7940 => state := s7941; 	--21
	addfpsclr <= '0';
when s7941 => state := s7942; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (416, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7942 => state := s7943; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (770, 12)); -- offset LSB 722
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s7943 => state := s7944;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (771, 12)); -- offset MSB 723
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7944 => state := s7945; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7945 => 			--4
	if (fixed2floatrdy = '1') then state := s7946;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7945; end if;
when s7946 => state := s7947; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7947 => 			--6
	if (mulfprdy = '1') then state := s7948;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7947; end if;
when s7948 => state := s7949; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7949 => 			--8
	if (mulfprdy = '1') then state := s7950;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7949; end if;
when s7950 => state := s7951; 	--9
	mulfpsclr <= '0';
when s7951 => state := s7952; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7952 => 			--11
	if (mulfprdy = '1') then state := s7953;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7952; end if;
when s7953 => state := s7954; 	--12
	mulfpsclr <= '0';
when s7954 => state := s7955; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7955 => 			--14
	if (addfprdy = '1') then state := s7956;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7955; end if;
when s7956 => state := s7957; 	--15
	addfpsclr <= '0';
when s7957 => state := s7958; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7958 => 			--17
	if (addfprdy = '1') then state := s7959;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7958; end if;
when s7959 => state := s7960; 	--18
	addfpsclr <= '0';
when s7960 => state := s7961; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7961 => 			--20
	if (addfprdy = '1') then state := s7962;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7961; end if;
when s7962 => state := s7963; 	--21
	addfpsclr <= '0';
when s7963 => state := s7964; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (417, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7964 => state := s7965; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (772, 12)); -- offset LSB 724
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s7965 => state := s7966;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (773, 12)); -- offset MSB 725
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7966 => state := s7967; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7967 => 			--4
	if (fixed2floatrdy = '1') then state := s7968;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7967; end if;
when s7968 => state := s7969; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7969 => 			--6
	if (mulfprdy = '1') then state := s7970;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7969; end if;
when s7970 => state := s7971; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7971 => 			--8
	if (mulfprdy = '1') then state := s7972;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7971; end if;
when s7972 => state := s7973; 	--9
	mulfpsclr <= '0';
when s7973 => state := s7974; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7974 => 			--11
	if (mulfprdy = '1') then state := s7975;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7974; end if;
when s7975 => state := s7976; 	--12
	mulfpsclr <= '0';
when s7976 => state := s7977; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7977 => 			--14
	if (addfprdy = '1') then state := s7978;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7977; end if;
when s7978 => state := s7979; 	--15
	addfpsclr <= '0';
when s7979 => state := s7980; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s7980 => 			--17
	if (addfprdy = '1') then state := s7981;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7980; end if;
when s7981 => state := s7982; 	--18
	addfpsclr <= '0';
when s7982 => state := s7983; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s7983 => 			--20
	if (addfprdy = '1') then state := s7984;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7983; end if;
when s7984 => state := s7985; 	--21
	addfpsclr <= '0';
when s7985 => state := s7986; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (418, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s7986 => state := s7987; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (774, 12)); -- offset LSB 726
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s7987 => state := s7988;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (775, 12)); -- offset MSB 727
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s7988 => state := s7989; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s7989 => 			--4
	if (fixed2floatrdy = '1') then state := s7990;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s7989; end if;
when s7990 => state := s7991; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s7991 => 			--6
	if (mulfprdy = '1') then state := s7992;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7991; end if;
when s7992 => state := s7993; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s7993 => 			--8
	if (mulfprdy = '1') then state := s7994;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7993; end if;
when s7994 => state := s7995; 	--9
	mulfpsclr <= '0';
when s7995 => state := s7996; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s7996 => 			--11
	if (mulfprdy = '1') then state := s7997;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s7996; end if;
when s7997 => state := s7998; 	--12
	mulfpsclr <= '0';
when s7998 => state := s7999; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s7999 => 			--14
	if (addfprdy = '1') then state := s8000;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s7999; end if;
when s8000 => state := s8001; 	--15
	addfpsclr <= '0';
when s8001 => state := s8002; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8002 => 			--17
	if (addfprdy = '1') then state := s8003;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8002; end if;
when s8003 => state := s8004; 	--18
	addfpsclr <= '0';
when s8004 => state := s8005; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8005 => 			--20
	if (addfprdy = '1') then state := s8006;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8005; end if;
when s8006 => state := s8007; 	--21
	addfpsclr <= '0';
when s8007 => state := s8008; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (419, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8008 => state := s8009; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (776, 12)); -- offset LSB 728
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s8009 => state := s8010;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (777, 12)); -- offset MSB 729
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8010 => state := s8011; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8011 => 			--4
	if (fixed2floatrdy = '1') then state := s8012;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8011; end if;
when s8012 => state := s8013; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8013 => 			--6
	if (mulfprdy = '1') then state := s8014;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8013; end if;
when s8014 => state := s8015; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8015 => 			--8
	if (mulfprdy = '1') then state := s8016;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8015; end if;
when s8016 => state := s8017; 	--9
	mulfpsclr <= '0';
when s8017 => state := s8018; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8018 => 			--11
	if (mulfprdy = '1') then state := s8019;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8018; end if;
when s8019 => state := s8020; 	--12
	mulfpsclr <= '0';
when s8020 => state := s8021; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8021 => 			--14
	if (addfprdy = '1') then state := s8022;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8021; end if;
when s8022 => state := s8023; 	--15
	addfpsclr <= '0';
when s8023 => state := s8024; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8024 => 			--17
	if (addfprdy = '1') then state := s8025;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8024; end if;
when s8025 => state := s8026; 	--18
	addfpsclr <= '0';
when s8026 => state := s8027; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8027 => 			--20
	if (addfprdy = '1') then state := s8028;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8027; end if;
when s8028 => state := s8029; 	--21
	addfpsclr <= '0';
when s8029 => state := s8030; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (420, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8030 => state := s8031; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (778, 12)); -- offset LSB 730
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s8031 => state := s8032;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (779, 12)); -- offset MSB 731
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8032 => state := s8033; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8033 => 			--4
	if (fixed2floatrdy = '1') then state := s8034;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8033; end if;
when s8034 => state := s8035; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8035 => 			--6
	if (mulfprdy = '1') then state := s8036;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8035; end if;
when s8036 => state := s8037; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8037 => 			--8
	if (mulfprdy = '1') then state := s8038;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8037; end if;
when s8038 => state := s8039; 	--9
	mulfpsclr <= '0';
when s8039 => state := s8040; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8040 => 			--11
	if (mulfprdy = '1') then state := s8041;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8040; end if;
when s8041 => state := s8042; 	--12
	mulfpsclr <= '0';
when s8042 => state := s8043; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8043 => 			--14
	if (addfprdy = '1') then state := s8044;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8043; end if;
when s8044 => state := s8045; 	--15
	addfpsclr <= '0';
when s8045 => state := s8046; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8046 => 			--17
	if (addfprdy = '1') then state := s8047;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8046; end if;
when s8047 => state := s8048; 	--18
	addfpsclr <= '0';
when s8048 => state := s8049; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8049 => 			--20
	if (addfprdy = '1') then state := s8050;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8049; end if;
when s8050 => state := s8051; 	--21
	addfpsclr <= '0';
when s8051 => state := s8052; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (421, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8052 => state := s8053; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (780, 12)); -- offset LSB 732
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s8053 => state := s8054;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (781, 12)); -- offset MSB 733
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8054 => state := s8055; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8055 => 			--4
	if (fixed2floatrdy = '1') then state := s8056;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8055; end if;
when s8056 => state := s8057; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8057 => 			--6
	if (mulfprdy = '1') then state := s8058;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8057; end if;
when s8058 => state := s8059; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8059 => 			--8
	if (mulfprdy = '1') then state := s8060;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8059; end if;
when s8060 => state := s8061; 	--9
	mulfpsclr <= '0';
when s8061 => state := s8062; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8062 => 			--11
	if (mulfprdy = '1') then state := s8063;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8062; end if;
when s8063 => state := s8064; 	--12
	mulfpsclr <= '0';
when s8064 => state := s8065; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8065 => 			--14
	if (addfprdy = '1') then state := s8066;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8065; end if;
when s8066 => state := s8067; 	--15
	addfpsclr <= '0';
when s8067 => state := s8068; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8068 => 			--17
	if (addfprdy = '1') then state := s8069;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8068; end if;
when s8069 => state := s8070; 	--18
	addfpsclr <= '0';
when s8070 => state := s8071; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8071 => 			--20
	if (addfprdy = '1') then state := s8072;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8071; end if;
when s8072 => state := s8073; 	--21
	addfpsclr <= '0';
when s8073 => state := s8074; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (422, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8074 => state := s8075; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (782, 12)); -- offset LSB 734
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s8075 => state := s8076;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (783, 12)); -- offset MSB 735
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8076 => state := s8077; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8077 => 			--4
	if (fixed2floatrdy = '1') then state := s8078;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8077; end if;
when s8078 => state := s8079; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8079 => 			--6
	if (mulfprdy = '1') then state := s8080;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8079; end if;
when s8080 => state := s8081; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8081 => 			--8
	if (mulfprdy = '1') then state := s8082;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8081; end if;
when s8082 => state := s8083; 	--9
	mulfpsclr <= '0';
when s8083 => state := s8084; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8084 => 			--11
	if (mulfprdy = '1') then state := s8085;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8084; end if;
when s8085 => state := s8086; 	--12
	mulfpsclr <= '0';
when s8086 => state := s8087; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8087 => 			--14
	if (addfprdy = '1') then state := s8088;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8087; end if;
when s8088 => state := s8089; 	--15
	addfpsclr <= '0';
when s8089 => state := s8090; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8090 => 			--17
	if (addfprdy = '1') then state := s8091;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8090; end if;
when s8091 => state := s8092; 	--18
	addfpsclr <= '0';
when s8092 => state := s8093; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8093 => 			--20
	if (addfprdy = '1') then state := s8094;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8093; end if;
when s8094 => state := s8095; 	--21
	addfpsclr <= '0';
when s8095 => state := s8096; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (423, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8096 => state := s8097; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (784, 12)); -- offset LSB 736
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s8097 => state := s8098;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (785, 12)); -- offset MSB 737
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8098 => state := s8099; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8099 => 			--4
	if (fixed2floatrdy = '1') then state := s8100;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8099; end if;
when s8100 => state := s8101; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8101 => 			--6
	if (mulfprdy = '1') then state := s8102;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8101; end if;
when s8102 => state := s8103; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8103 => 			--8
	if (mulfprdy = '1') then state := s8104;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8103; end if;
when s8104 => state := s8105; 	--9
	mulfpsclr <= '0';
when s8105 => state := s8106; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8106 => 			--11
	if (mulfprdy = '1') then state := s8107;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8106; end if;
when s8107 => state := s8108; 	--12
	mulfpsclr <= '0';
when s8108 => state := s8109; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8109 => 			--14
	if (addfprdy = '1') then state := s8110;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8109; end if;
when s8110 => state := s8111; 	--15
	addfpsclr <= '0';
when s8111 => state := s8112; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8112 => 			--17
	if (addfprdy = '1') then state := s8113;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8112; end if;
when s8113 => state := s8114; 	--18
	addfpsclr <= '0';
when s8114 => state := s8115; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8115 => 			--20
	if (addfprdy = '1') then state := s8116;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8115; end if;
when s8116 => state := s8117; 	--21
	addfpsclr <= '0';
when s8117 => state := s8118; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (424, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8118 => state := s8119; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (786, 12)); -- offset LSB 738
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s8119 => state := s8120;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (787, 12)); -- offset MSB 739
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8120 => state := s8121; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8121 => 			--4
	if (fixed2floatrdy = '1') then state := s8122;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8121; end if;
when s8122 => state := s8123; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8123 => 			--6
	if (mulfprdy = '1') then state := s8124;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8123; end if;
when s8124 => state := s8125; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8125 => 			--8
	if (mulfprdy = '1') then state := s8126;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8125; end if;
when s8126 => state := s8127; 	--9
	mulfpsclr <= '0';
when s8127 => state := s8128; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8128 => 			--11
	if (mulfprdy = '1') then state := s8129;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8128; end if;
when s8129 => state := s8130; 	--12
	mulfpsclr <= '0';
when s8130 => state := s8131; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8131 => 			--14
	if (addfprdy = '1') then state := s8132;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8131; end if;
when s8132 => state := s8133; 	--15
	addfpsclr <= '0';
when s8133 => state := s8134; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8134 => 			--17
	if (addfprdy = '1') then state := s8135;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8134; end if;
when s8135 => state := s8136; 	--18
	addfpsclr <= '0';
when s8136 => state := s8137; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8137 => 			--20
	if (addfprdy = '1') then state := s8138;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8137; end if;
when s8138 => state := s8139; 	--21
	addfpsclr <= '0';
when s8139 => state := s8140; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (425, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8140 => state := s8141; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (788, 12)); -- offset LSB 740
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s8141 => state := s8142;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (789, 12)); -- offset MSB 741
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8142 => state := s8143; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8143 => 			--4
	if (fixed2floatrdy = '1') then state := s8144;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8143; end if;
when s8144 => state := s8145; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8145 => 			--6
	if (mulfprdy = '1') then state := s8146;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8145; end if;
when s8146 => state := s8147; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8147 => 			--8
	if (mulfprdy = '1') then state := s8148;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8147; end if;
when s8148 => state := s8149; 	--9
	mulfpsclr <= '0';
when s8149 => state := s8150; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8150 => 			--11
	if (mulfprdy = '1') then state := s8151;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8150; end if;
when s8151 => state := s8152; 	--12
	mulfpsclr <= '0';
when s8152 => state := s8153; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8153 => 			--14
	if (addfprdy = '1') then state := s8154;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8153; end if;
when s8154 => state := s8155; 	--15
	addfpsclr <= '0';
when s8155 => state := s8156; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8156 => 			--17
	if (addfprdy = '1') then state := s8157;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8156; end if;
when s8157 => state := s8158; 	--18
	addfpsclr <= '0';
when s8158 => state := s8159; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8159 => 			--20
	if (addfprdy = '1') then state := s8160;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8159; end if;
when s8160 => state := s8161; 	--21
	addfpsclr <= '0';
when s8161 => state := s8162; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (426, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8162 => state := s8163; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (790, 12)); -- offset LSB 742
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s8163 => state := s8164;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (791, 12)); -- offset MSB 743
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8164 => state := s8165; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8165 => 			--4
	if (fixed2floatrdy = '1') then state := s8166;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8165; end if;
when s8166 => state := s8167; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8167 => 			--6
	if (mulfprdy = '1') then state := s8168;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8167; end if;
when s8168 => state := s8169; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8169 => 			--8
	if (mulfprdy = '1') then state := s8170;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8169; end if;
when s8170 => state := s8171; 	--9
	mulfpsclr <= '0';
when s8171 => state := s8172; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8172 => 			--11
	if (mulfprdy = '1') then state := s8173;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8172; end if;
when s8173 => state := s8174; 	--12
	mulfpsclr <= '0';
when s8174 => state := s8175; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8175 => 			--14
	if (addfprdy = '1') then state := s8176;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8175; end if;
when s8176 => state := s8177; 	--15
	addfpsclr <= '0';
when s8177 => state := s8178; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8178 => 			--17
	if (addfprdy = '1') then state := s8179;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8178; end if;
when s8179 => state := s8180; 	--18
	addfpsclr <= '0';
when s8180 => state := s8181; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8181 => 			--20
	if (addfprdy = '1') then state := s8182;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8181; end if;
when s8182 => state := s8183; 	--21
	addfpsclr <= '0';
when s8183 => state := s8184; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (427, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8184 => state := s8185; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (792, 12)); -- offset LSB 744
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s8185 => state := s8186;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (793, 12)); -- offset MSB 745
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8186 => state := s8187; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8187 => 			--4
	if (fixed2floatrdy = '1') then state := s8188;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8187; end if;
when s8188 => state := s8189; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8189 => 			--6
	if (mulfprdy = '1') then state := s8190;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8189; end if;
when s8190 => state := s8191; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8191 => 			--8
	if (mulfprdy = '1') then state := s8192;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8191; end if;
when s8192 => state := s8193; 	--9
	mulfpsclr <= '0';
when s8193 => state := s8194; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8194 => 			--11
	if (mulfprdy = '1') then state := s8195;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8194; end if;
when s8195 => state := s8196; 	--12
	mulfpsclr <= '0';
when s8196 => state := s8197; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8197 => 			--14
	if (addfprdy = '1') then state := s8198;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8197; end if;
when s8198 => state := s8199; 	--15
	addfpsclr <= '0';
when s8199 => state := s8200; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8200 => 			--17
	if (addfprdy = '1') then state := s8201;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8200; end if;
when s8201 => state := s8202; 	--18
	addfpsclr <= '0';
when s8202 => state := s8203; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8203 => 			--20
	if (addfprdy = '1') then state := s8204;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8203; end if;
when s8204 => state := s8205; 	--21
	addfpsclr <= '0';
when s8205 => state := s8206; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (428, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8206 => state := s8207; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (794, 12)); -- offset LSB 746
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s8207 => state := s8208;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (795, 12)); -- offset MSB 747
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8208 => state := s8209; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8209 => 			--4
	if (fixed2floatrdy = '1') then state := s8210;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8209; end if;
when s8210 => state := s8211; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8211 => 			--6
	if (mulfprdy = '1') then state := s8212;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8211; end if;
when s8212 => state := s8213; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8213 => 			--8
	if (mulfprdy = '1') then state := s8214;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8213; end if;
when s8214 => state := s8215; 	--9
	mulfpsclr <= '0';
when s8215 => state := s8216; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8216 => 			--11
	if (mulfprdy = '1') then state := s8217;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8216; end if;
when s8217 => state := s8218; 	--12
	mulfpsclr <= '0';
when s8218 => state := s8219; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8219 => 			--14
	if (addfprdy = '1') then state := s8220;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8219; end if;
when s8220 => state := s8221; 	--15
	addfpsclr <= '0';
when s8221 => state := s8222; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8222 => 			--17
	if (addfprdy = '1') then state := s8223;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8222; end if;
when s8223 => state := s8224; 	--18
	addfpsclr <= '0';
when s8224 => state := s8225; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8225 => 			--20
	if (addfprdy = '1') then state := s8226;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8225; end if;
when s8226 => state := s8227; 	--21
	addfpsclr <= '0';
when s8227 => state := s8228; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (429, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8228 => state := s8229; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (796, 12)); -- offset LSB 748
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s8229 => state := s8230;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (797, 12)); -- offset MSB 749
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8230 => state := s8231; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8231 => 			--4
	if (fixed2floatrdy = '1') then state := s8232;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8231; end if;
when s8232 => state := s8233; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8233 => 			--6
	if (mulfprdy = '1') then state := s8234;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8233; end if;
when s8234 => state := s8235; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8235 => 			--8
	if (mulfprdy = '1') then state := s8236;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8235; end if;
when s8236 => state := s8237; 	--9
	mulfpsclr <= '0';
when s8237 => state := s8238; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8238 => 			--11
	if (mulfprdy = '1') then state := s8239;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8238; end if;
when s8239 => state := s8240; 	--12
	mulfpsclr <= '0';
when s8240 => state := s8241; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8241 => 			--14
	if (addfprdy = '1') then state := s8242;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8241; end if;
when s8242 => state := s8243; 	--15
	addfpsclr <= '0';
when s8243 => state := s8244; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8244 => 			--17
	if (addfprdy = '1') then state := s8245;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8244; end if;
when s8245 => state := s8246; 	--18
	addfpsclr <= '0';
when s8246 => state := s8247; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8247 => 			--20
	if (addfprdy = '1') then state := s8248;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8247; end if;
when s8248 => state := s8249; 	--21
	addfpsclr <= '0';
when s8249 => state := s8250; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (430, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8250 => state := s8251; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (798, 12)); -- offset LSB 750
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s8251 => state := s8252;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (799, 12)); -- offset MSB 751
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8252 => state := s8253; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8253 => 			--4
	if (fixed2floatrdy = '1') then state := s8254;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8253; end if;
when s8254 => state := s8255; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8255 => 			--6
	if (mulfprdy = '1') then state := s8256;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8255; end if;
when s8256 => state := s8257; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8257 => 			--8
	if (mulfprdy = '1') then state := s8258;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8257; end if;
when s8258 => state := s8259; 	--9
	mulfpsclr <= '0';
when s8259 => state := s8260; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8260 => 			--11
	if (mulfprdy = '1') then state := s8261;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8260; end if;
when s8261 => state := s8262; 	--12
	mulfpsclr <= '0';
when s8262 => state := s8263; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8263 => 			--14
	if (addfprdy = '1') then state := s8264;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8263; end if;
when s8264 => state := s8265; 	--15
	addfpsclr <= '0';
when s8265 => state := s8266; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8266 => 			--17
	if (addfprdy = '1') then state := s8267;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8266; end if;
when s8267 => state := s8268; 	--18
	addfpsclr <= '0';
when s8268 => state := s8269; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8269 => 			--20
	if (addfprdy = '1') then state := s8270;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8269; end if;
when s8270 => state := s8271; 	--21
	addfpsclr <= '0';
when s8271 => state := s8272; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (431, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8272 => state := s8273; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (800, 12)); -- offset LSB 752
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s8273 => state := s8274;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (801, 12)); -- offset MSB 753
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8274 => state := s8275; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8275 => 			--4
	if (fixed2floatrdy = '1') then state := s8276;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8275; end if;
when s8276 => state := s8277; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8277 => 			--6
	if (mulfprdy = '1') then state := s8278;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8277; end if;
when s8278 => state := s8279; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8279 => 			--8
	if (mulfprdy = '1') then state := s8280;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8279; end if;
when s8280 => state := s8281; 	--9
	mulfpsclr <= '0';
when s8281 => state := s8282; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8282 => 			--11
	if (mulfprdy = '1') then state := s8283;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8282; end if;
when s8283 => state := s8284; 	--12
	mulfpsclr <= '0';
when s8284 => state := s8285; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8285 => 			--14
	if (addfprdy = '1') then state := s8286;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8285; end if;
when s8286 => state := s8287; 	--15
	addfpsclr <= '0';
when s8287 => state := s8288; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8288 => 			--17
	if (addfprdy = '1') then state := s8289;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8288; end if;
when s8289 => state := s8290; 	--18
	addfpsclr <= '0';
when s8290 => state := s8291; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8291 => 			--20
	if (addfprdy = '1') then state := s8292;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8291; end if;
when s8292 => state := s8293; 	--21
	addfpsclr <= '0';
when s8293 => state := s8294; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (432, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8294 => state := s8295; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (802, 12)); -- offset LSB 754
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s8295 => state := s8296;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (803, 12)); -- offset MSB 755
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8296 => state := s8297; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8297 => 			--4
	if (fixed2floatrdy = '1') then state := s8298;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8297; end if;
when s8298 => state := s8299; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8299 => 			--6
	if (mulfprdy = '1') then state := s8300;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8299; end if;
when s8300 => state := s8301; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8301 => 			--8
	if (mulfprdy = '1') then state := s8302;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8301; end if;
when s8302 => state := s8303; 	--9
	mulfpsclr <= '0';
when s8303 => state := s8304; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8304 => 			--11
	if (mulfprdy = '1') then state := s8305;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8304; end if;
when s8305 => state := s8306; 	--12
	mulfpsclr <= '0';
when s8306 => state := s8307; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8307 => 			--14
	if (addfprdy = '1') then state := s8308;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8307; end if;
when s8308 => state := s8309; 	--15
	addfpsclr <= '0';
when s8309 => state := s8310; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8310 => 			--17
	if (addfprdy = '1') then state := s8311;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8310; end if;
when s8311 => state := s8312; 	--18
	addfpsclr <= '0';
when s8312 => state := s8313; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8313 => 			--20
	if (addfprdy = '1') then state := s8314;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8313; end if;
when s8314 => state := s8315; 	--21
	addfpsclr <= '0';
when s8315 => state := s8316; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (433, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8316 => state := s8317; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (804, 12)); -- offset LSB 756
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s8317 => state := s8318;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (805, 12)); -- offset MSB 757
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8318 => state := s8319; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8319 => 			--4
	if (fixed2floatrdy = '1') then state := s8320;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8319; end if;
when s8320 => state := s8321; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8321 => 			--6
	if (mulfprdy = '1') then state := s8322;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8321; end if;
when s8322 => state := s8323; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8323 => 			--8
	if (mulfprdy = '1') then state := s8324;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8323; end if;
when s8324 => state := s8325; 	--9
	mulfpsclr <= '0';
when s8325 => state := s8326; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8326 => 			--11
	if (mulfprdy = '1') then state := s8327;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8326; end if;
when s8327 => state := s8328; 	--12
	mulfpsclr <= '0';
when s8328 => state := s8329; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8329 => 			--14
	if (addfprdy = '1') then state := s8330;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8329; end if;
when s8330 => state := s8331; 	--15
	addfpsclr <= '0';
when s8331 => state := s8332; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8332 => 			--17
	if (addfprdy = '1') then state := s8333;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8332; end if;
when s8333 => state := s8334; 	--18
	addfpsclr <= '0';
when s8334 => state := s8335; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8335 => 			--20
	if (addfprdy = '1') then state := s8336;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8335; end if;
when s8336 => state := s8337; 	--21
	addfpsclr <= '0';
when s8337 => state := s8338; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (434, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8338 => state := s8339; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (806, 12)); -- offset LSB 758
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s8339 => state := s8340;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (807, 12)); -- offset MSB 759
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8340 => state := s8341; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8341 => 			--4
	if (fixed2floatrdy = '1') then state := s8342;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8341; end if;
when s8342 => state := s8343; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8343 => 			--6
	if (mulfprdy = '1') then state := s8344;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8343; end if;
when s8344 => state := s8345; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8345 => 			--8
	if (mulfprdy = '1') then state := s8346;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8345; end if;
when s8346 => state := s8347; 	--9
	mulfpsclr <= '0';
when s8347 => state := s8348; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8348 => 			--11
	if (mulfprdy = '1') then state := s8349;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8348; end if;
when s8349 => state := s8350; 	--12
	mulfpsclr <= '0';
when s8350 => state := s8351; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8351 => 			--14
	if (addfprdy = '1') then state := s8352;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8351; end if;
when s8352 => state := s8353; 	--15
	addfpsclr <= '0';
when s8353 => state := s8354; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8354 => 			--17
	if (addfprdy = '1') then state := s8355;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8354; end if;
when s8355 => state := s8356; 	--18
	addfpsclr <= '0';
when s8356 => state := s8357; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8357 => 			--20
	if (addfprdy = '1') then state := s8358;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8357; end if;
when s8358 => state := s8359; 	--21
	addfpsclr <= '0';
when s8359 => state := s8360; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (435, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8360 => state := s8361; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (808, 12)); -- offset LSB 760
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s8361 => state := s8362;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (809, 12)); -- offset MSB 761
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8362 => state := s8363; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8363 => 			--4
	if (fixed2floatrdy = '1') then state := s8364;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8363; end if;
when s8364 => state := s8365; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8365 => 			--6
	if (mulfprdy = '1') then state := s8366;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8365; end if;
when s8366 => state := s8367; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8367 => 			--8
	if (mulfprdy = '1') then state := s8368;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8367; end if;
when s8368 => state := s8369; 	--9
	mulfpsclr <= '0';
when s8369 => state := s8370; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8370 => 			--11
	if (mulfprdy = '1') then state := s8371;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8370; end if;
when s8371 => state := s8372; 	--12
	mulfpsclr <= '0';
when s8372 => state := s8373; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8373 => 			--14
	if (addfprdy = '1') then state := s8374;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8373; end if;
when s8374 => state := s8375; 	--15
	addfpsclr <= '0';
when s8375 => state := s8376; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8376 => 			--17
	if (addfprdy = '1') then state := s8377;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8376; end if;
when s8377 => state := s8378; 	--18
	addfpsclr <= '0';
when s8378 => state := s8379; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8379 => 			--20
	if (addfprdy = '1') then state := s8380;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8379; end if;
when s8380 => state := s8381; 	--21
	addfpsclr <= '0';
when s8381 => state := s8382; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (436, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8382 => state := s8383; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (810, 12)); -- offset LSB 762
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s8383 => state := s8384;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (811, 12)); -- offset MSB 763
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8384 => state := s8385; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8385 => 			--4
	if (fixed2floatrdy = '1') then state := s8386;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8385; end if;
when s8386 => state := s8387; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8387 => 			--6
	if (mulfprdy = '1') then state := s8388;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8387; end if;
when s8388 => state := s8389; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8389 => 			--8
	if (mulfprdy = '1') then state := s8390;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8389; end if;
when s8390 => state := s8391; 	--9
	mulfpsclr <= '0';
when s8391 => state := s8392; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8392 => 			--11
	if (mulfprdy = '1') then state := s8393;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8392; end if;
when s8393 => state := s8394; 	--12
	mulfpsclr <= '0';
when s8394 => state := s8395; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8395 => 			--14
	if (addfprdy = '1') then state := s8396;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8395; end if;
when s8396 => state := s8397; 	--15
	addfpsclr <= '0';
when s8397 => state := s8398; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8398 => 			--17
	if (addfprdy = '1') then state := s8399;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8398; end if;
when s8399 => state := s8400; 	--18
	addfpsclr <= '0';
when s8400 => state := s8401; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8401 => 			--20
	if (addfprdy = '1') then state := s8402;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8401; end if;
when s8402 => state := s8403; 	--21
	addfpsclr <= '0';
when s8403 => state := s8404; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (437, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8404 => state := s8405; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (812, 12)); -- offset LSB 764
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s8405 => state := s8406;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (813, 12)); -- offset MSB 765
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8406 => state := s8407; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8407 => 			--4
	if (fixed2floatrdy = '1') then state := s8408;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8407; end if;
when s8408 => state := s8409; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8409 => 			--6
	if (mulfprdy = '1') then state := s8410;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8409; end if;
when s8410 => state := s8411; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8411 => 			--8
	if (mulfprdy = '1') then state := s8412;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8411; end if;
when s8412 => state := s8413; 	--9
	mulfpsclr <= '0';
when s8413 => state := s8414; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8414 => 			--11
	if (mulfprdy = '1') then state := s8415;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8414; end if;
when s8415 => state := s8416; 	--12
	mulfpsclr <= '0';
when s8416 => state := s8417; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8417 => 			--14
	if (addfprdy = '1') then state := s8418;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8417; end if;
when s8418 => state := s8419; 	--15
	addfpsclr <= '0';
when s8419 => state := s8420; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8420 => 			--17
	if (addfprdy = '1') then state := s8421;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8420; end if;
when s8421 => state := s8422; 	--18
	addfpsclr <= '0';
when s8422 => state := s8423; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8423 => 			--20
	if (addfprdy = '1') then state := s8424;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8423; end if;
when s8424 => state := s8425; 	--21
	addfpsclr <= '0';
when s8425 => state := s8426; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (438, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8426 => state := s8427; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (814, 12)); -- offset LSB 766
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s8427 => state := s8428;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (815, 12)); -- offset MSB 767
	addra <= std_logic_vector (to_unsigned (11, 10)); -- OCCrowI 11
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8428 => state := s8429; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8429 => 			--4
	if (fixed2floatrdy = '1') then state := s8430;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8429; end if;
when s8430 => state := s8431; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8431 => 			--6
	if (mulfprdy = '1') then state := s8432;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8431; end if;
when s8432 => state := s8433; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8433 => 			--8
	if (mulfprdy = '1') then state := s8434;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8433; end if;
when s8434 => state := s8435; 	--9
	mulfpsclr <= '0';
when s8435 => state := s8436; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8436 => 			--11
	if (mulfprdy = '1') then state := s8437;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8436; end if;
when s8437 => state := s8438; 	--12
	mulfpsclr <= '0';
when s8438 => state := s8439; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8439 => 			--14
	if (addfprdy = '1') then state := s8440;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8439; end if;
when s8440 => state := s8441; 	--15
	addfpsclr <= '0';
when s8441 => state := s8442; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8442 => 			--17
	if (addfprdy = '1') then state := s8443;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8442; end if;
when s8443 => state := s8444; 	--18
	addfpsclr <= '0';
when s8444 => state := s8445; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8445 => 			--20
	if (addfprdy = '1') then state := s8446;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8445; end if;
when s8446 => state := s8447; 	--21
	addfpsclr <= '0';
when s8447 => state := s8448; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (439, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8448 => state := s8449; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (816, 12)); -- offset LSB 768
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s8449 => state := s8450;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (817, 12)); -- offset MSB 769
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8450 => state := s8451; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8451 => 			--4
	if (fixed2floatrdy = '1') then state := s8452;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8451; end if;
when s8452 => state := s8453; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8453 => 			--6
	if (mulfprdy = '1') then state := s8454;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8453; end if;
when s8454 => state := s8455; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8455 => 			--8
	if (mulfprdy = '1') then state := s8456;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8455; end if;
when s8456 => state := s8457; 	--9
	mulfpsclr <= '0';
when s8457 => state := s8458; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8458 => 			--11
	if (mulfprdy = '1') then state := s8459;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8458; end if;
when s8459 => state := s8460; 	--12
	mulfpsclr <= '0';
when s8460 => state := s8461; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8461 => 			--14
	if (addfprdy = '1') then state := s8462;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8461; end if;
when s8462 => state := s8463; 	--15
	addfpsclr <= '0';
when s8463 => state := s8464; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8464 => 			--17
	if (addfprdy = '1') then state := s8465;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8464; end if;
when s8465 => state := s8466; 	--18
	addfpsclr <= '0';
when s8466 => state := s8467; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8467 => 			--20
	if (addfprdy = '1') then state := s8468;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8467; end if;
when s8468 => state := s8469; 	--21
	addfpsclr <= '0';
when s8469 => state := s8470; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (440, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8470 => state := s8471; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (818, 12)); -- offset LSB 770
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s8471 => state := s8472;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (819, 12)); -- offset MSB 771
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8472 => state := s8473; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8473 => 			--4
	if (fixed2floatrdy = '1') then state := s8474;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8473; end if;
when s8474 => state := s8475; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8475 => 			--6
	if (mulfprdy = '1') then state := s8476;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8475; end if;
when s8476 => state := s8477; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8477 => 			--8
	if (mulfprdy = '1') then state := s8478;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8477; end if;
when s8478 => state := s8479; 	--9
	mulfpsclr <= '0';
when s8479 => state := s8480; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8480 => 			--11
	if (mulfprdy = '1') then state := s8481;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8480; end if;
when s8481 => state := s8482; 	--12
	mulfpsclr <= '0';
when s8482 => state := s8483; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8483 => 			--14
	if (addfprdy = '1') then state := s8484;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8483; end if;
when s8484 => state := s8485; 	--15
	addfpsclr <= '0';
when s8485 => state := s8486; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8486 => 			--17
	if (addfprdy = '1') then state := s8487;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8486; end if;
when s8487 => state := s8488; 	--18
	addfpsclr <= '0';
when s8488 => state := s8489; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8489 => 			--20
	if (addfprdy = '1') then state := s8490;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8489; end if;
when s8490 => state := s8491; 	--21
	addfpsclr <= '0';
when s8491 => state := s8492; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (441, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8492 => state := s8493; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (820, 12)); -- offset LSB 772
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s8493 => state := s8494;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (821, 12)); -- offset MSB 773
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8494 => state := s8495; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8495 => 			--4
	if (fixed2floatrdy = '1') then state := s8496;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8495; end if;
when s8496 => state := s8497; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8497 => 			--6
	if (mulfprdy = '1') then state := s8498;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8497; end if;
when s8498 => state := s8499; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8499 => 			--8
	if (mulfprdy = '1') then state := s8500;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8499; end if;
when s8500 => state := s8501; 	--9
	mulfpsclr <= '0';
when s8501 => state := s8502; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8502 => 			--11
	if (mulfprdy = '1') then state := s8503;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8502; end if;
when s8503 => state := s8504; 	--12
	mulfpsclr <= '0';
when s8504 => state := s8505; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8505 => 			--14
	if (addfprdy = '1') then state := s8506;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8505; end if;
when s8506 => state := s8507; 	--15
	addfpsclr <= '0';
when s8507 => state := s8508; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8508 => 			--17
	if (addfprdy = '1') then state := s8509;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8508; end if;
when s8509 => state := s8510; 	--18
	addfpsclr <= '0';
when s8510 => state := s8511; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8511 => 			--20
	if (addfprdy = '1') then state := s8512;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8511; end if;
when s8512 => state := s8513; 	--21
	addfpsclr <= '0';
when s8513 => state := s8514; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (442, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8514 => state := s8515; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (822, 12)); -- offset LSB 774
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s8515 => state := s8516;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (823, 12)); -- offset MSB 775
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8516 => state := s8517; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8517 => 			--4
	if (fixed2floatrdy = '1') then state := s8518;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8517; end if;
when s8518 => state := s8519; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8519 => 			--6
	if (mulfprdy = '1') then state := s8520;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8519; end if;
when s8520 => state := s8521; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8521 => 			--8
	if (mulfprdy = '1') then state := s8522;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8521; end if;
when s8522 => state := s8523; 	--9
	mulfpsclr <= '0';
when s8523 => state := s8524; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8524 => 			--11
	if (mulfprdy = '1') then state := s8525;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8524; end if;
when s8525 => state := s8526; 	--12
	mulfpsclr <= '0';
when s8526 => state := s8527; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8527 => 			--14
	if (addfprdy = '1') then state := s8528;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8527; end if;
when s8528 => state := s8529; 	--15
	addfpsclr <= '0';
when s8529 => state := s8530; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8530 => 			--17
	if (addfprdy = '1') then state := s8531;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8530; end if;
when s8531 => state := s8532; 	--18
	addfpsclr <= '0';
when s8532 => state := s8533; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8533 => 			--20
	if (addfprdy = '1') then state := s8534;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8533; end if;
when s8534 => state := s8535; 	--21
	addfpsclr <= '0';
when s8535 => state := s8536; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (443, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8536 => state := s8537; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (824, 12)); -- offset LSB 776
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s8537 => state := s8538;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (825, 12)); -- offset MSB 777
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8538 => state := s8539; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8539 => 			--4
	if (fixed2floatrdy = '1') then state := s8540;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8539; end if;
when s8540 => state := s8541; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8541 => 			--6
	if (mulfprdy = '1') then state := s8542;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8541; end if;
when s8542 => state := s8543; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8543 => 			--8
	if (mulfprdy = '1') then state := s8544;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8543; end if;
when s8544 => state := s8545; 	--9
	mulfpsclr <= '0';
when s8545 => state := s8546; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8546 => 			--11
	if (mulfprdy = '1') then state := s8547;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8546; end if;
when s8547 => state := s8548; 	--12
	mulfpsclr <= '0';
when s8548 => state := s8549; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8549 => 			--14
	if (addfprdy = '1') then state := s8550;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8549; end if;
when s8550 => state := s8551; 	--15
	addfpsclr <= '0';
when s8551 => state := s8552; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8552 => 			--17
	if (addfprdy = '1') then state := s8553;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8552; end if;
when s8553 => state := s8554; 	--18
	addfpsclr <= '0';
when s8554 => state := s8555; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8555 => 			--20
	if (addfprdy = '1') then state := s8556;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8555; end if;
when s8556 => state := s8557; 	--21
	addfpsclr <= '0';
when s8557 => state := s8558; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (444, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8558 => state := s8559; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (826, 12)); -- offset LSB 778
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s8559 => state := s8560;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (827, 12)); -- offset MSB 779
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8560 => state := s8561; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8561 => 			--4
	if (fixed2floatrdy = '1') then state := s8562;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8561; end if;
when s8562 => state := s8563; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8563 => 			--6
	if (mulfprdy = '1') then state := s8564;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8563; end if;
when s8564 => state := s8565; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8565 => 			--8
	if (mulfprdy = '1') then state := s8566;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8565; end if;
when s8566 => state := s8567; 	--9
	mulfpsclr <= '0';
when s8567 => state := s8568; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8568 => 			--11
	if (mulfprdy = '1') then state := s8569;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8568; end if;
when s8569 => state := s8570; 	--12
	mulfpsclr <= '0';
when s8570 => state := s8571; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8571 => 			--14
	if (addfprdy = '1') then state := s8572;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8571; end if;
when s8572 => state := s8573; 	--15
	addfpsclr <= '0';
when s8573 => state := s8574; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8574 => 			--17
	if (addfprdy = '1') then state := s8575;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8574; end if;
when s8575 => state := s8576; 	--18
	addfpsclr <= '0';
when s8576 => state := s8577; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8577 => 			--20
	if (addfprdy = '1') then state := s8578;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8577; end if;
when s8578 => state := s8579; 	--21
	addfpsclr <= '0';
when s8579 => state := s8580; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (445, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8580 => state := s8581; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (828, 12)); -- offset LSB 780
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s8581 => state := s8582;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (829, 12)); -- offset MSB 781
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8582 => state := s8583; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8583 => 			--4
	if (fixed2floatrdy = '1') then state := s8584;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8583; end if;
when s8584 => state := s8585; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8585 => 			--6
	if (mulfprdy = '1') then state := s8586;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8585; end if;
when s8586 => state := s8587; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8587 => 			--8
	if (mulfprdy = '1') then state := s8588;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8587; end if;
when s8588 => state := s8589; 	--9
	mulfpsclr <= '0';
when s8589 => state := s8590; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8590 => 			--11
	if (mulfprdy = '1') then state := s8591;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8590; end if;
when s8591 => state := s8592; 	--12
	mulfpsclr <= '0';
when s8592 => state := s8593; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8593 => 			--14
	if (addfprdy = '1') then state := s8594;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8593; end if;
when s8594 => state := s8595; 	--15
	addfpsclr <= '0';
when s8595 => state := s8596; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8596 => 			--17
	if (addfprdy = '1') then state := s8597;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8596; end if;
when s8597 => state := s8598; 	--18
	addfpsclr <= '0';
when s8598 => state := s8599; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8599 => 			--20
	if (addfprdy = '1') then state := s8600;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8599; end if;
when s8600 => state := s8601; 	--21
	addfpsclr <= '0';
when s8601 => state := s8602; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (446, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8602 => state := s8603; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (830, 12)); -- offset LSB 782
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s8603 => state := s8604;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (831, 12)); -- offset MSB 783
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8604 => state := s8605; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8605 => 			--4
	if (fixed2floatrdy = '1') then state := s8606;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8605; end if;
when s8606 => state := s8607; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8607 => 			--6
	if (mulfprdy = '1') then state := s8608;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8607; end if;
when s8608 => state := s8609; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8609 => 			--8
	if (mulfprdy = '1') then state := s8610;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8609; end if;
when s8610 => state := s8611; 	--9
	mulfpsclr <= '0';
when s8611 => state := s8612; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8612 => 			--11
	if (mulfprdy = '1') then state := s8613;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8612; end if;
when s8613 => state := s8614; 	--12
	mulfpsclr <= '0';
when s8614 => state := s8615; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8615 => 			--14
	if (addfprdy = '1') then state := s8616;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8615; end if;
when s8616 => state := s8617; 	--15
	addfpsclr <= '0';
when s8617 => state := s8618; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8618 => 			--17
	if (addfprdy = '1') then state := s8619;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8618; end if;
when s8619 => state := s8620; 	--18
	addfpsclr <= '0';
when s8620 => state := s8621; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8621 => 			--20
	if (addfprdy = '1') then state := s8622;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8621; end if;
when s8622 => state := s8623; 	--21
	addfpsclr <= '0';
when s8623 => state := s8624; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (447, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8624 => state := s8625; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (832, 12)); -- offset LSB 784
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s8625 => state := s8626;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (833, 12)); -- offset MSB 785
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8626 => state := s8627; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8627 => 			--4
	if (fixed2floatrdy = '1') then state := s8628;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8627; end if;
when s8628 => state := s8629; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8629 => 			--6
	if (mulfprdy = '1') then state := s8630;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8629; end if;
when s8630 => state := s8631; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8631 => 			--8
	if (mulfprdy = '1') then state := s8632;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8631; end if;
when s8632 => state := s8633; 	--9
	mulfpsclr <= '0';
when s8633 => state := s8634; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8634 => 			--11
	if (mulfprdy = '1') then state := s8635;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8634; end if;
when s8635 => state := s8636; 	--12
	mulfpsclr <= '0';
when s8636 => state := s8637; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8637 => 			--14
	if (addfprdy = '1') then state := s8638;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8637; end if;
when s8638 => state := s8639; 	--15
	addfpsclr <= '0';
when s8639 => state := s8640; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8640 => 			--17
	if (addfprdy = '1') then state := s8641;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8640; end if;
when s8641 => state := s8642; 	--18
	addfpsclr <= '0';
when s8642 => state := s8643; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8643 => 			--20
	if (addfprdy = '1') then state := s8644;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8643; end if;
when s8644 => state := s8645; 	--21
	addfpsclr <= '0';
when s8645 => state := s8646; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (448, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8646 => state := s8647; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (834, 12)); -- offset LSB 786
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s8647 => state := s8648;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (835, 12)); -- offset MSB 787
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8648 => state := s8649; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8649 => 			--4
	if (fixed2floatrdy = '1') then state := s8650;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8649; end if;
when s8650 => state := s8651; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8651 => 			--6
	if (mulfprdy = '1') then state := s8652;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8651; end if;
when s8652 => state := s8653; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8653 => 			--8
	if (mulfprdy = '1') then state := s8654;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8653; end if;
when s8654 => state := s8655; 	--9
	mulfpsclr <= '0';
when s8655 => state := s8656; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8656 => 			--11
	if (mulfprdy = '1') then state := s8657;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8656; end if;
when s8657 => state := s8658; 	--12
	mulfpsclr <= '0';
when s8658 => state := s8659; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8659 => 			--14
	if (addfprdy = '1') then state := s8660;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8659; end if;
when s8660 => state := s8661; 	--15
	addfpsclr <= '0';
when s8661 => state := s8662; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8662 => 			--17
	if (addfprdy = '1') then state := s8663;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8662; end if;
when s8663 => state := s8664; 	--18
	addfpsclr <= '0';
when s8664 => state := s8665; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8665 => 			--20
	if (addfprdy = '1') then state := s8666;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8665; end if;
when s8666 => state := s8667; 	--21
	addfpsclr <= '0';
when s8667 => state := s8668; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (449, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8668 => state := s8669; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (836, 12)); -- offset LSB 788
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s8669 => state := s8670;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (837, 12)); -- offset MSB 789
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8670 => state := s8671; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8671 => 			--4
	if (fixed2floatrdy = '1') then state := s8672;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8671; end if;
when s8672 => state := s8673; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8673 => 			--6
	if (mulfprdy = '1') then state := s8674;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8673; end if;
when s8674 => state := s8675; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8675 => 			--8
	if (mulfprdy = '1') then state := s8676;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8675; end if;
when s8676 => state := s8677; 	--9
	mulfpsclr <= '0';
when s8677 => state := s8678; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8678 => 			--11
	if (mulfprdy = '1') then state := s8679;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8678; end if;
when s8679 => state := s8680; 	--12
	mulfpsclr <= '0';
when s8680 => state := s8681; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8681 => 			--14
	if (addfprdy = '1') then state := s8682;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8681; end if;
when s8682 => state := s8683; 	--15
	addfpsclr <= '0';
when s8683 => state := s8684; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8684 => 			--17
	if (addfprdy = '1') then state := s8685;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8684; end if;
when s8685 => state := s8686; 	--18
	addfpsclr <= '0';
when s8686 => state := s8687; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8687 => 			--20
	if (addfprdy = '1') then state := s8688;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8687; end if;
when s8688 => state := s8689; 	--21
	addfpsclr <= '0';
when s8689 => state := s8690; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (450, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8690 => state := s8691; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (838, 12)); -- offset LSB 790
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s8691 => state := s8692;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (839, 12)); -- offset MSB 791
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8692 => state := s8693; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8693 => 			--4
	if (fixed2floatrdy = '1') then state := s8694;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8693; end if;
when s8694 => state := s8695; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8695 => 			--6
	if (mulfprdy = '1') then state := s8696;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8695; end if;
when s8696 => state := s8697; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8697 => 			--8
	if (mulfprdy = '1') then state := s8698;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8697; end if;
when s8698 => state := s8699; 	--9
	mulfpsclr <= '0';
when s8699 => state := s8700; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8700 => 			--11
	if (mulfprdy = '1') then state := s8701;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8700; end if;
when s8701 => state := s8702; 	--12
	mulfpsclr <= '0';
when s8702 => state := s8703; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8703 => 			--14
	if (addfprdy = '1') then state := s8704;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8703; end if;
when s8704 => state := s8705; 	--15
	addfpsclr <= '0';
when s8705 => state := s8706; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8706 => 			--17
	if (addfprdy = '1') then state := s8707;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8706; end if;
when s8707 => state := s8708; 	--18
	addfpsclr <= '0';
when s8708 => state := s8709; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8709 => 			--20
	if (addfprdy = '1') then state := s8710;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8709; end if;
when s8710 => state := s8711; 	--21
	addfpsclr <= '0';
when s8711 => state := s8712; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (451, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8712 => state := s8713; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (840, 12)); -- offset LSB 792
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s8713 => state := s8714;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (841, 12)); -- offset MSB 793
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8714 => state := s8715; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8715 => 			--4
	if (fixed2floatrdy = '1') then state := s8716;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8715; end if;
when s8716 => state := s8717; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8717 => 			--6
	if (mulfprdy = '1') then state := s8718;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8717; end if;
when s8718 => state := s8719; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8719 => 			--8
	if (mulfprdy = '1') then state := s8720;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8719; end if;
when s8720 => state := s8721; 	--9
	mulfpsclr <= '0';
when s8721 => state := s8722; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8722 => 			--11
	if (mulfprdy = '1') then state := s8723;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8722; end if;
when s8723 => state := s8724; 	--12
	mulfpsclr <= '0';
when s8724 => state := s8725; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8725 => 			--14
	if (addfprdy = '1') then state := s8726;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8725; end if;
when s8726 => state := s8727; 	--15
	addfpsclr <= '0';
when s8727 => state := s8728; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8728 => 			--17
	if (addfprdy = '1') then state := s8729;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8728; end if;
when s8729 => state := s8730; 	--18
	addfpsclr <= '0';
when s8730 => state := s8731; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8731 => 			--20
	if (addfprdy = '1') then state := s8732;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8731; end if;
when s8732 => state := s8733; 	--21
	addfpsclr <= '0';
when s8733 => state := s8734; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (452, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8734 => state := s8735; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (842, 12)); -- offset LSB 794
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s8735 => state := s8736;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (843, 12)); -- offset MSB 795
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8736 => state := s8737; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8737 => 			--4
	if (fixed2floatrdy = '1') then state := s8738;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8737; end if;
when s8738 => state := s8739; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8739 => 			--6
	if (mulfprdy = '1') then state := s8740;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8739; end if;
when s8740 => state := s8741; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8741 => 			--8
	if (mulfprdy = '1') then state := s8742;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8741; end if;
when s8742 => state := s8743; 	--9
	mulfpsclr <= '0';
when s8743 => state := s8744; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8744 => 			--11
	if (mulfprdy = '1') then state := s8745;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8744; end if;
when s8745 => state := s8746; 	--12
	mulfpsclr <= '0';
when s8746 => state := s8747; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8747 => 			--14
	if (addfprdy = '1') then state := s8748;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8747; end if;
when s8748 => state := s8749; 	--15
	addfpsclr <= '0';
when s8749 => state := s8750; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8750 => 			--17
	if (addfprdy = '1') then state := s8751;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8750; end if;
when s8751 => state := s8752; 	--18
	addfpsclr <= '0';
when s8752 => state := s8753; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8753 => 			--20
	if (addfprdy = '1') then state := s8754;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8753; end if;
when s8754 => state := s8755; 	--21
	addfpsclr <= '0';
when s8755 => state := s8756; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (453, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8756 => state := s8757; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (844, 12)); -- offset LSB 796
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s8757 => state := s8758;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (845, 12)); -- offset MSB 797
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8758 => state := s8759; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8759 => 			--4
	if (fixed2floatrdy = '1') then state := s8760;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8759; end if;
when s8760 => state := s8761; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8761 => 			--6
	if (mulfprdy = '1') then state := s8762;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8761; end if;
when s8762 => state := s8763; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8763 => 			--8
	if (mulfprdy = '1') then state := s8764;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8763; end if;
when s8764 => state := s8765; 	--9
	mulfpsclr <= '0';
when s8765 => state := s8766; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8766 => 			--11
	if (mulfprdy = '1') then state := s8767;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8766; end if;
when s8767 => state := s8768; 	--12
	mulfpsclr <= '0';
when s8768 => state := s8769; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8769 => 			--14
	if (addfprdy = '1') then state := s8770;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8769; end if;
when s8770 => state := s8771; 	--15
	addfpsclr <= '0';
when s8771 => state := s8772; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8772 => 			--17
	if (addfprdy = '1') then state := s8773;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8772; end if;
when s8773 => state := s8774; 	--18
	addfpsclr <= '0';
when s8774 => state := s8775; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8775 => 			--20
	if (addfprdy = '1') then state := s8776;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8775; end if;
when s8776 => state := s8777; 	--21
	addfpsclr <= '0';
when s8777 => state := s8778; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (454, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8778 => state := s8779; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (846, 12)); -- offset LSB 798
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s8779 => state := s8780;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (847, 12)); -- offset MSB 799
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8780 => state := s8781; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8781 => 			--4
	if (fixed2floatrdy = '1') then state := s8782;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8781; end if;
when s8782 => state := s8783; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8783 => 			--6
	if (mulfprdy = '1') then state := s8784;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8783; end if;
when s8784 => state := s8785; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8785 => 			--8
	if (mulfprdy = '1') then state := s8786;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8785; end if;
when s8786 => state := s8787; 	--9
	mulfpsclr <= '0';
when s8787 => state := s8788; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8788 => 			--11
	if (mulfprdy = '1') then state := s8789;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8788; end if;
when s8789 => state := s8790; 	--12
	mulfpsclr <= '0';
when s8790 => state := s8791; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8791 => 			--14
	if (addfprdy = '1') then state := s8792;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8791; end if;
when s8792 => state := s8793; 	--15
	addfpsclr <= '0';
when s8793 => state := s8794; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8794 => 			--17
	if (addfprdy = '1') then state := s8795;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8794; end if;
when s8795 => state := s8796; 	--18
	addfpsclr <= '0';
when s8796 => state := s8797; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8797 => 			--20
	if (addfprdy = '1') then state := s8798;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8797; end if;
when s8798 => state := s8799; 	--21
	addfpsclr <= '0';
when s8799 => state := s8800; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (455, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8800 => state := s8801; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (848, 12)); -- offset LSB 800
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s8801 => state := s8802;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (849, 12)); -- offset MSB 801
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8802 => state := s8803; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8803 => 			--4
	if (fixed2floatrdy = '1') then state := s8804;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8803; end if;
when s8804 => state := s8805; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8805 => 			--6
	if (mulfprdy = '1') then state := s8806;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8805; end if;
when s8806 => state := s8807; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8807 => 			--8
	if (mulfprdy = '1') then state := s8808;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8807; end if;
when s8808 => state := s8809; 	--9
	mulfpsclr <= '0';
when s8809 => state := s8810; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8810 => 			--11
	if (mulfprdy = '1') then state := s8811;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8810; end if;
when s8811 => state := s8812; 	--12
	mulfpsclr <= '0';
when s8812 => state := s8813; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8813 => 			--14
	if (addfprdy = '1') then state := s8814;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8813; end if;
when s8814 => state := s8815; 	--15
	addfpsclr <= '0';
when s8815 => state := s8816; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8816 => 			--17
	if (addfprdy = '1') then state := s8817;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8816; end if;
when s8817 => state := s8818; 	--18
	addfpsclr <= '0';
when s8818 => state := s8819; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8819 => 			--20
	if (addfprdy = '1') then state := s8820;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8819; end if;
when s8820 => state := s8821; 	--21
	addfpsclr <= '0';
when s8821 => state := s8822; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (456, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8822 => state := s8823; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (850, 12)); -- offset LSB 802
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s8823 => state := s8824;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (851, 12)); -- offset MSB 803
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8824 => state := s8825; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8825 => 			--4
	if (fixed2floatrdy = '1') then state := s8826;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8825; end if;
when s8826 => state := s8827; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8827 => 			--6
	if (mulfprdy = '1') then state := s8828;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8827; end if;
when s8828 => state := s8829; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8829 => 			--8
	if (mulfprdy = '1') then state := s8830;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8829; end if;
when s8830 => state := s8831; 	--9
	mulfpsclr <= '0';
when s8831 => state := s8832; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8832 => 			--11
	if (mulfprdy = '1') then state := s8833;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8832; end if;
when s8833 => state := s8834; 	--12
	mulfpsclr <= '0';
when s8834 => state := s8835; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8835 => 			--14
	if (addfprdy = '1') then state := s8836;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8835; end if;
when s8836 => state := s8837; 	--15
	addfpsclr <= '0';
when s8837 => state := s8838; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8838 => 			--17
	if (addfprdy = '1') then state := s8839;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8838; end if;
when s8839 => state := s8840; 	--18
	addfpsclr <= '0';
when s8840 => state := s8841; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8841 => 			--20
	if (addfprdy = '1') then state := s8842;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8841; end if;
when s8842 => state := s8843; 	--21
	addfpsclr <= '0';
when s8843 => state := s8844; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (457, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8844 => state := s8845; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (852, 12)); -- offset LSB 804
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s8845 => state := s8846;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (853, 12)); -- offset MSB 805
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8846 => state := s8847; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8847 => 			--4
	if (fixed2floatrdy = '1') then state := s8848;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8847; end if;
when s8848 => state := s8849; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8849 => 			--6
	if (mulfprdy = '1') then state := s8850;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8849; end if;
when s8850 => state := s8851; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8851 => 			--8
	if (mulfprdy = '1') then state := s8852;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8851; end if;
when s8852 => state := s8853; 	--9
	mulfpsclr <= '0';
when s8853 => state := s8854; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8854 => 			--11
	if (mulfprdy = '1') then state := s8855;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8854; end if;
when s8855 => state := s8856; 	--12
	mulfpsclr <= '0';
when s8856 => state := s8857; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8857 => 			--14
	if (addfprdy = '1') then state := s8858;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8857; end if;
when s8858 => state := s8859; 	--15
	addfpsclr <= '0';
when s8859 => state := s8860; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8860 => 			--17
	if (addfprdy = '1') then state := s8861;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8860; end if;
when s8861 => state := s8862; 	--18
	addfpsclr <= '0';
when s8862 => state := s8863; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8863 => 			--20
	if (addfprdy = '1') then state := s8864;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8863; end if;
when s8864 => state := s8865; 	--21
	addfpsclr <= '0';
when s8865 => state := s8866; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (458, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8866 => state := s8867; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (854, 12)); -- offset LSB 806
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s8867 => state := s8868;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (855, 12)); -- offset MSB 807
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8868 => state := s8869; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8869 => 			--4
	if (fixed2floatrdy = '1') then state := s8870;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8869; end if;
when s8870 => state := s8871; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8871 => 			--6
	if (mulfprdy = '1') then state := s8872;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8871; end if;
when s8872 => state := s8873; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8873 => 			--8
	if (mulfprdy = '1') then state := s8874;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8873; end if;
when s8874 => state := s8875; 	--9
	mulfpsclr <= '0';
when s8875 => state := s8876; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8876 => 			--11
	if (mulfprdy = '1') then state := s8877;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8876; end if;
when s8877 => state := s8878; 	--12
	mulfpsclr <= '0';
when s8878 => state := s8879; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8879 => 			--14
	if (addfprdy = '1') then state := s8880;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8879; end if;
when s8880 => state := s8881; 	--15
	addfpsclr <= '0';
when s8881 => state := s8882; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8882 => 			--17
	if (addfprdy = '1') then state := s8883;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8882; end if;
when s8883 => state := s8884; 	--18
	addfpsclr <= '0';
when s8884 => state := s8885; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8885 => 			--20
	if (addfprdy = '1') then state := s8886;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8885; end if;
when s8886 => state := s8887; 	--21
	addfpsclr <= '0';
when s8887 => state := s8888; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (459, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8888 => state := s8889; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (856, 12)); -- offset LSB 808
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s8889 => state := s8890;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (857, 12)); -- offset MSB 809
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8890 => state := s8891; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8891 => 			--4
	if (fixed2floatrdy = '1') then state := s8892;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8891; end if;
when s8892 => state := s8893; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8893 => 			--6
	if (mulfprdy = '1') then state := s8894;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8893; end if;
when s8894 => state := s8895; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8895 => 			--8
	if (mulfprdy = '1') then state := s8896;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8895; end if;
when s8896 => state := s8897; 	--9
	mulfpsclr <= '0';
when s8897 => state := s8898; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8898 => 			--11
	if (mulfprdy = '1') then state := s8899;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8898; end if;
when s8899 => state := s8900; 	--12
	mulfpsclr <= '0';
when s8900 => state := s8901; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8901 => 			--14
	if (addfprdy = '1') then state := s8902;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8901; end if;
when s8902 => state := s8903; 	--15
	addfpsclr <= '0';
when s8903 => state := s8904; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8904 => 			--17
	if (addfprdy = '1') then state := s8905;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8904; end if;
when s8905 => state := s8906; 	--18
	addfpsclr <= '0';
when s8906 => state := s8907; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8907 => 			--20
	if (addfprdy = '1') then state := s8908;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8907; end if;
when s8908 => state := s8909; 	--21
	addfpsclr <= '0';
when s8909 => state := s8910; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (460, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8910 => state := s8911; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (858, 12)); -- offset LSB 810
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s8911 => state := s8912;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (859, 12)); -- offset MSB 811
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8912 => state := s8913; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8913 => 			--4
	if (fixed2floatrdy = '1') then state := s8914;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8913; end if;
when s8914 => state := s8915; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8915 => 			--6
	if (mulfprdy = '1') then state := s8916;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8915; end if;
when s8916 => state := s8917; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8917 => 			--8
	if (mulfprdy = '1') then state := s8918;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8917; end if;
when s8918 => state := s8919; 	--9
	mulfpsclr <= '0';
when s8919 => state := s8920; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8920 => 			--11
	if (mulfprdy = '1') then state := s8921;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8920; end if;
when s8921 => state := s8922; 	--12
	mulfpsclr <= '0';
when s8922 => state := s8923; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8923 => 			--14
	if (addfprdy = '1') then state := s8924;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8923; end if;
when s8924 => state := s8925; 	--15
	addfpsclr <= '0';
when s8925 => state := s8926; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8926 => 			--17
	if (addfprdy = '1') then state := s8927;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8926; end if;
when s8927 => state := s8928; 	--18
	addfpsclr <= '0';
when s8928 => state := s8929; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8929 => 			--20
	if (addfprdy = '1') then state := s8930;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8929; end if;
when s8930 => state := s8931; 	--21
	addfpsclr <= '0';
when s8931 => state := s8932; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (461, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8932 => state := s8933; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (860, 12)); -- offset LSB 812
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s8933 => state := s8934;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (861, 12)); -- offset MSB 813
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8934 => state := s8935; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8935 => 			--4
	if (fixed2floatrdy = '1') then state := s8936;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8935; end if;
when s8936 => state := s8937; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8937 => 			--6
	if (mulfprdy = '1') then state := s8938;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8937; end if;
when s8938 => state := s8939; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8939 => 			--8
	if (mulfprdy = '1') then state := s8940;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8939; end if;
when s8940 => state := s8941; 	--9
	mulfpsclr <= '0';
when s8941 => state := s8942; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8942 => 			--11
	if (mulfprdy = '1') then state := s8943;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8942; end if;
when s8943 => state := s8944; 	--12
	mulfpsclr <= '0';
when s8944 => state := s8945; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8945 => 			--14
	if (addfprdy = '1') then state := s8946;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8945; end if;
when s8946 => state := s8947; 	--15
	addfpsclr <= '0';
when s8947 => state := s8948; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8948 => 			--17
	if (addfprdy = '1') then state := s8949;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8948; end if;
when s8949 => state := s8950; 	--18
	addfpsclr <= '0';
when s8950 => state := s8951; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8951 => 			--20
	if (addfprdy = '1') then state := s8952;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8951; end if;
when s8952 => state := s8953; 	--21
	addfpsclr <= '0';
when s8953 => state := s8954; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (462, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8954 => state := s8955; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (862, 12)); -- offset LSB 814
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s8955 => state := s8956;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (863, 12)); -- offset MSB 815
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8956 => state := s8957; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8957 => 			--4
	if (fixed2floatrdy = '1') then state := s8958;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8957; end if;
when s8958 => state := s8959; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8959 => 			--6
	if (mulfprdy = '1') then state := s8960;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8959; end if;
when s8960 => state := s8961; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8961 => 			--8
	if (mulfprdy = '1') then state := s8962;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8961; end if;
when s8962 => state := s8963; 	--9
	mulfpsclr <= '0';
when s8963 => state := s8964; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8964 => 			--11
	if (mulfprdy = '1') then state := s8965;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8964; end if;
when s8965 => state := s8966; 	--12
	mulfpsclr <= '0';
when s8966 => state := s8967; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8967 => 			--14
	if (addfprdy = '1') then state := s8968;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8967; end if;
when s8968 => state := s8969; 	--15
	addfpsclr <= '0';
when s8969 => state := s8970; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8970 => 			--17
	if (addfprdy = '1') then state := s8971;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8970; end if;
when s8971 => state := s8972; 	--18
	addfpsclr <= '0';
when s8972 => state := s8973; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8973 => 			--20
	if (addfprdy = '1') then state := s8974;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8973; end if;
when s8974 => state := s8975; 	--21
	addfpsclr <= '0';
when s8975 => state := s8976; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (463, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8976 => state := s8977; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (864, 12)); -- offset LSB 816
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s8977 => state := s8978;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (865, 12)); -- offset MSB 817
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s8978 => state := s8979; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s8979 => 			--4
	if (fixed2floatrdy = '1') then state := s8980;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s8979; end if;
when s8980 => state := s8981; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s8981 => 			--6
	if (mulfprdy = '1') then state := s8982;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8981; end if;
when s8982 => state := s8983; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s8983 => 			--8
	if (mulfprdy = '1') then state := s8984;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8983; end if;
when s8984 => state := s8985; 	--9
	mulfpsclr <= '0';
when s8985 => state := s8986; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s8986 => 			--11
	if (mulfprdy = '1') then state := s8987;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s8986; end if;
when s8987 => state := s8988; 	--12
	mulfpsclr <= '0';
when s8988 => state := s8989; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s8989 => 			--14
	if (addfprdy = '1') then state := s8990;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8989; end if;
when s8990 => state := s8991; 	--15
	addfpsclr <= '0';
when s8991 => state := s8992; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s8992 => 			--17
	if (addfprdy = '1') then state := s8993;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8992; end if;
when s8993 => state := s8994; 	--18
	addfpsclr <= '0';
when s8994 => state := s8995; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s8995 => 			--20
	if (addfprdy = '1') then state := s8996;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s8995; end if;
when s8996 => state := s8997; 	--21
	addfpsclr <= '0';
when s8997 => state := s8998; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (464, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s8998 => state := s8999; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (866, 12)); -- offset LSB 818
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s8999 => state := s9000;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (867, 12)); -- offset MSB 819
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9000 => state := s9001; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9001 => 			--4
	if (fixed2floatrdy = '1') then state := s9002;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9001; end if;
when s9002 => state := s9003; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9003 => 			--6
	if (mulfprdy = '1') then state := s9004;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9003; end if;
when s9004 => state := s9005; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9005 => 			--8
	if (mulfprdy = '1') then state := s9006;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9005; end if;
when s9006 => state := s9007; 	--9
	mulfpsclr <= '0';
when s9007 => state := s9008; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9008 => 			--11
	if (mulfprdy = '1') then state := s9009;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9008; end if;
when s9009 => state := s9010; 	--12
	mulfpsclr <= '0';
when s9010 => state := s9011; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9011 => 			--14
	if (addfprdy = '1') then state := s9012;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9011; end if;
when s9012 => state := s9013; 	--15
	addfpsclr <= '0';
when s9013 => state := s9014; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9014 => 			--17
	if (addfprdy = '1') then state := s9015;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9014; end if;
when s9015 => state := s9016; 	--18
	addfpsclr <= '0';
when s9016 => state := s9017; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9017 => 			--20
	if (addfprdy = '1') then state := s9018;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9017; end if;
when s9018 => state := s9019; 	--21
	addfpsclr <= '0';
when s9019 => state := s9020; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (465, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9020 => state := s9021; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (868, 12)); -- offset LSB 820
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s9021 => state := s9022;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (869, 12)); -- offset MSB 821
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9022 => state := s9023; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9023 => 			--4
	if (fixed2floatrdy = '1') then state := s9024;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9023; end if;
when s9024 => state := s9025; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9025 => 			--6
	if (mulfprdy = '1') then state := s9026;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9025; end if;
when s9026 => state := s9027; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9027 => 			--8
	if (mulfprdy = '1') then state := s9028;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9027; end if;
when s9028 => state := s9029; 	--9
	mulfpsclr <= '0';
when s9029 => state := s9030; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9030 => 			--11
	if (mulfprdy = '1') then state := s9031;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9030; end if;
when s9031 => state := s9032; 	--12
	mulfpsclr <= '0';
when s9032 => state := s9033; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9033 => 			--14
	if (addfprdy = '1') then state := s9034;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9033; end if;
when s9034 => state := s9035; 	--15
	addfpsclr <= '0';
when s9035 => state := s9036; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9036 => 			--17
	if (addfprdy = '1') then state := s9037;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9036; end if;
when s9037 => state := s9038; 	--18
	addfpsclr <= '0';
when s9038 => state := s9039; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9039 => 			--20
	if (addfprdy = '1') then state := s9040;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9039; end if;
when s9040 => state := s9041; 	--21
	addfpsclr <= '0';
when s9041 => state := s9042; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (466, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9042 => state := s9043; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (870, 12)); -- offset LSB 822
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s9043 => state := s9044;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (871, 12)); -- offset MSB 823
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9044 => state := s9045; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9045 => 			--4
	if (fixed2floatrdy = '1') then state := s9046;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9045; end if;
when s9046 => state := s9047; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9047 => 			--6
	if (mulfprdy = '1') then state := s9048;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9047; end if;
when s9048 => state := s9049; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9049 => 			--8
	if (mulfprdy = '1') then state := s9050;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9049; end if;
when s9050 => state := s9051; 	--9
	mulfpsclr <= '0';
when s9051 => state := s9052; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9052 => 			--11
	if (mulfprdy = '1') then state := s9053;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9052; end if;
when s9053 => state := s9054; 	--12
	mulfpsclr <= '0';
when s9054 => state := s9055; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9055 => 			--14
	if (addfprdy = '1') then state := s9056;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9055; end if;
when s9056 => state := s9057; 	--15
	addfpsclr <= '0';
when s9057 => state := s9058; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9058 => 			--17
	if (addfprdy = '1') then state := s9059;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9058; end if;
when s9059 => state := s9060; 	--18
	addfpsclr <= '0';
when s9060 => state := s9061; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9061 => 			--20
	if (addfprdy = '1') then state := s9062;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9061; end if;
when s9062 => state := s9063; 	--21
	addfpsclr <= '0';
when s9063 => state := s9064; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (467, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9064 => state := s9065; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (872, 12)); -- offset LSB 824
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s9065 => state := s9066;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (873, 12)); -- offset MSB 825
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9066 => state := s9067; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9067 => 			--4
	if (fixed2floatrdy = '1') then state := s9068;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9067; end if;
when s9068 => state := s9069; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9069 => 			--6
	if (mulfprdy = '1') then state := s9070;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9069; end if;
when s9070 => state := s9071; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9071 => 			--8
	if (mulfprdy = '1') then state := s9072;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9071; end if;
when s9072 => state := s9073; 	--9
	mulfpsclr <= '0';
when s9073 => state := s9074; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9074 => 			--11
	if (mulfprdy = '1') then state := s9075;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9074; end if;
when s9075 => state := s9076; 	--12
	mulfpsclr <= '0';
when s9076 => state := s9077; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9077 => 			--14
	if (addfprdy = '1') then state := s9078;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9077; end if;
when s9078 => state := s9079; 	--15
	addfpsclr <= '0';
when s9079 => state := s9080; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9080 => 			--17
	if (addfprdy = '1') then state := s9081;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9080; end if;
when s9081 => state := s9082; 	--18
	addfpsclr <= '0';
when s9082 => state := s9083; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9083 => 			--20
	if (addfprdy = '1') then state := s9084;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9083; end if;
when s9084 => state := s9085; 	--21
	addfpsclr <= '0';
when s9085 => state := s9086; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (468, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9086 => state := s9087; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (874, 12)); -- offset LSB 826
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s9087 => state := s9088;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (875, 12)); -- offset MSB 827
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9088 => state := s9089; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9089 => 			--4
	if (fixed2floatrdy = '1') then state := s9090;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9089; end if;
when s9090 => state := s9091; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9091 => 			--6
	if (mulfprdy = '1') then state := s9092;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9091; end if;
when s9092 => state := s9093; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9093 => 			--8
	if (mulfprdy = '1') then state := s9094;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9093; end if;
when s9094 => state := s9095; 	--9
	mulfpsclr <= '0';
when s9095 => state := s9096; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9096 => 			--11
	if (mulfprdy = '1') then state := s9097;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9096; end if;
when s9097 => state := s9098; 	--12
	mulfpsclr <= '0';
when s9098 => state := s9099; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9099 => 			--14
	if (addfprdy = '1') then state := s9100;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9099; end if;
when s9100 => state := s9101; 	--15
	addfpsclr <= '0';
when s9101 => state := s9102; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9102 => 			--17
	if (addfprdy = '1') then state := s9103;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9102; end if;
when s9103 => state := s9104; 	--18
	addfpsclr <= '0';
when s9104 => state := s9105; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9105 => 			--20
	if (addfprdy = '1') then state := s9106;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9105; end if;
when s9106 => state := s9107; 	--21
	addfpsclr <= '0';
when s9107 => state := s9108; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (469, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9108 => state := s9109; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (876, 12)); -- offset LSB 828
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s9109 => state := s9110;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (877, 12)); -- offset MSB 829
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9110 => state := s9111; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9111 => 			--4
	if (fixed2floatrdy = '1') then state := s9112;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9111; end if;
when s9112 => state := s9113; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9113 => 			--6
	if (mulfprdy = '1') then state := s9114;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9113; end if;
when s9114 => state := s9115; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9115 => 			--8
	if (mulfprdy = '1') then state := s9116;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9115; end if;
when s9116 => state := s9117; 	--9
	mulfpsclr <= '0';
when s9117 => state := s9118; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9118 => 			--11
	if (mulfprdy = '1') then state := s9119;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9118; end if;
when s9119 => state := s9120; 	--12
	mulfpsclr <= '0';
when s9120 => state := s9121; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9121 => 			--14
	if (addfprdy = '1') then state := s9122;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9121; end if;
when s9122 => state := s9123; 	--15
	addfpsclr <= '0';
when s9123 => state := s9124; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9124 => 			--17
	if (addfprdy = '1') then state := s9125;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9124; end if;
when s9125 => state := s9126; 	--18
	addfpsclr <= '0';
when s9126 => state := s9127; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9127 => 			--20
	if (addfprdy = '1') then state := s9128;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9127; end if;
when s9128 => state := s9129; 	--21
	addfpsclr <= '0';
when s9129 => state := s9130; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (470, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9130 => state := s9131; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (878, 12)); -- offset LSB 830
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s9131 => state := s9132;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (879, 12)); -- offset MSB 831
	addra <= std_logic_vector (to_unsigned (12, 10)); -- OCCrowI 12
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9132 => state := s9133; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9133 => 			--4
	if (fixed2floatrdy = '1') then state := s9134;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9133; end if;
when s9134 => state := s9135; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9135 => 			--6
	if (mulfprdy = '1') then state := s9136;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9135; end if;
when s9136 => state := s9137; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9137 => 			--8
	if (mulfprdy = '1') then state := s9138;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9137; end if;
when s9138 => state := s9139; 	--9
	mulfpsclr <= '0';
when s9139 => state := s9140; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9140 => 			--11
	if (mulfprdy = '1') then state := s9141;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9140; end if;
when s9141 => state := s9142; 	--12
	mulfpsclr <= '0';
when s9142 => state := s9143; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9143 => 			--14
	if (addfprdy = '1') then state := s9144;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9143; end if;
when s9144 => state := s9145; 	--15
	addfpsclr <= '0';
when s9145 => state := s9146; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9146 => 			--17
	if (addfprdy = '1') then state := s9147;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9146; end if;
when s9147 => state := s9148; 	--18
	addfpsclr <= '0';
when s9148 => state := s9149; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9149 => 			--20
	if (addfprdy = '1') then state := s9150;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9149; end if;
when s9150 => state := s9151; 	--21
	addfpsclr <= '0';
when s9151 => state := s9152; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (471, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9152 => state := s9153; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (880, 12)); -- offset LSB 832
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s9153 => state := s9154;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (881, 12)); -- offset MSB 833
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9154 => state := s9155; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9155 => 			--4
	if (fixed2floatrdy = '1') then state := s9156;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9155; end if;
when s9156 => state := s9157; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9157 => 			--6
	if (mulfprdy = '1') then state := s9158;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9157; end if;
when s9158 => state := s9159; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9159 => 			--8
	if (mulfprdy = '1') then state := s9160;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9159; end if;
when s9160 => state := s9161; 	--9
	mulfpsclr <= '0';
when s9161 => state := s9162; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9162 => 			--11
	if (mulfprdy = '1') then state := s9163;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9162; end if;
when s9163 => state := s9164; 	--12
	mulfpsclr <= '0';
when s9164 => state := s9165; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9165 => 			--14
	if (addfprdy = '1') then state := s9166;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9165; end if;
when s9166 => state := s9167; 	--15
	addfpsclr <= '0';
when s9167 => state := s9168; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9168 => 			--17
	if (addfprdy = '1') then state := s9169;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9168; end if;
when s9169 => state := s9170; 	--18
	addfpsclr <= '0';
when s9170 => state := s9171; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9171 => 			--20
	if (addfprdy = '1') then state := s9172;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9171; end if;
when s9172 => state := s9173; 	--21
	addfpsclr <= '0';
when s9173 => state := s9174; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (472, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9174 => state := s9175; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (882, 12)); -- offset LSB 834
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s9175 => state := s9176;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (883, 12)); -- offset MSB 835
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9176 => state := s9177; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9177 => 			--4
	if (fixed2floatrdy = '1') then state := s9178;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9177; end if;
when s9178 => state := s9179; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9179 => 			--6
	if (mulfprdy = '1') then state := s9180;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9179; end if;
when s9180 => state := s9181; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9181 => 			--8
	if (mulfprdy = '1') then state := s9182;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9181; end if;
when s9182 => state := s9183; 	--9
	mulfpsclr <= '0';
when s9183 => state := s9184; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9184 => 			--11
	if (mulfprdy = '1') then state := s9185;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9184; end if;
when s9185 => state := s9186; 	--12
	mulfpsclr <= '0';
when s9186 => state := s9187; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9187 => 			--14
	if (addfprdy = '1') then state := s9188;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9187; end if;
when s9188 => state := s9189; 	--15
	addfpsclr <= '0';
when s9189 => state := s9190; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9190 => 			--17
	if (addfprdy = '1') then state := s9191;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9190; end if;
when s9191 => state := s9192; 	--18
	addfpsclr <= '0';
when s9192 => state := s9193; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9193 => 			--20
	if (addfprdy = '1') then state := s9194;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9193; end if;
when s9194 => state := s9195; 	--21
	addfpsclr <= '0';
when s9195 => state := s9196; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (473, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9196 => state := s9197; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (884, 12)); -- offset LSB 836
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s9197 => state := s9198;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (885, 12)); -- offset MSB 837
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9198 => state := s9199; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9199 => 			--4
	if (fixed2floatrdy = '1') then state := s9200;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9199; end if;
when s9200 => state := s9201; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9201 => 			--6
	if (mulfprdy = '1') then state := s9202;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9201; end if;
when s9202 => state := s9203; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9203 => 			--8
	if (mulfprdy = '1') then state := s9204;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9203; end if;
when s9204 => state := s9205; 	--9
	mulfpsclr <= '0';
when s9205 => state := s9206; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9206 => 			--11
	if (mulfprdy = '1') then state := s9207;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9206; end if;
when s9207 => state := s9208; 	--12
	mulfpsclr <= '0';
when s9208 => state := s9209; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9209 => 			--14
	if (addfprdy = '1') then state := s9210;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9209; end if;
when s9210 => state := s9211; 	--15
	addfpsclr <= '0';
when s9211 => state := s9212; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9212 => 			--17
	if (addfprdy = '1') then state := s9213;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9212; end if;
when s9213 => state := s9214; 	--18
	addfpsclr <= '0';
when s9214 => state := s9215; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9215 => 			--20
	if (addfprdy = '1') then state := s9216;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9215; end if;
when s9216 => state := s9217; 	--21
	addfpsclr <= '0';
when s9217 => state := s9218; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (474, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9218 => state := s9219; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (886, 12)); -- offset LSB 838
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s9219 => state := s9220;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (887, 12)); -- offset MSB 839
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9220 => state := s9221; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9221 => 			--4
	if (fixed2floatrdy = '1') then state := s9222;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9221; end if;
when s9222 => state := s9223; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9223 => 			--6
	if (mulfprdy = '1') then state := s9224;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9223; end if;
when s9224 => state := s9225; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9225 => 			--8
	if (mulfprdy = '1') then state := s9226;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9225; end if;
when s9226 => state := s9227; 	--9
	mulfpsclr <= '0';
when s9227 => state := s9228; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9228 => 			--11
	if (mulfprdy = '1') then state := s9229;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9228; end if;
when s9229 => state := s9230; 	--12
	mulfpsclr <= '0';
when s9230 => state := s9231; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9231 => 			--14
	if (addfprdy = '1') then state := s9232;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9231; end if;
when s9232 => state := s9233; 	--15
	addfpsclr <= '0';
when s9233 => state := s9234; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9234 => 			--17
	if (addfprdy = '1') then state := s9235;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9234; end if;
when s9235 => state := s9236; 	--18
	addfpsclr <= '0';
when s9236 => state := s9237; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9237 => 			--20
	if (addfprdy = '1') then state := s9238;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9237; end if;
when s9238 => state := s9239; 	--21
	addfpsclr <= '0';
when s9239 => state := s9240; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (475, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9240 => state := s9241; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (888, 12)); -- offset LSB 840
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s9241 => state := s9242;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (889, 12)); -- offset MSB 841
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9242 => state := s9243; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9243 => 			--4
	if (fixed2floatrdy = '1') then state := s9244;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9243; end if;
when s9244 => state := s9245; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9245 => 			--6
	if (mulfprdy = '1') then state := s9246;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9245; end if;
when s9246 => state := s9247; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9247 => 			--8
	if (mulfprdy = '1') then state := s9248;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9247; end if;
when s9248 => state := s9249; 	--9
	mulfpsclr <= '0';
when s9249 => state := s9250; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9250 => 			--11
	if (mulfprdy = '1') then state := s9251;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9250; end if;
when s9251 => state := s9252; 	--12
	mulfpsclr <= '0';
when s9252 => state := s9253; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9253 => 			--14
	if (addfprdy = '1') then state := s9254;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9253; end if;
when s9254 => state := s9255; 	--15
	addfpsclr <= '0';
when s9255 => state := s9256; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9256 => 			--17
	if (addfprdy = '1') then state := s9257;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9256; end if;
when s9257 => state := s9258; 	--18
	addfpsclr <= '0';
when s9258 => state := s9259; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9259 => 			--20
	if (addfprdy = '1') then state := s9260;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9259; end if;
when s9260 => state := s9261; 	--21
	addfpsclr <= '0';
when s9261 => state := s9262; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (476, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9262 => state := s9263; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (890, 12)); -- offset LSB 842
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s9263 => state := s9264;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (891, 12)); -- offset MSB 843
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9264 => state := s9265; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9265 => 			--4
	if (fixed2floatrdy = '1') then state := s9266;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9265; end if;
when s9266 => state := s9267; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9267 => 			--6
	if (mulfprdy = '1') then state := s9268;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9267; end if;
when s9268 => state := s9269; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9269 => 			--8
	if (mulfprdy = '1') then state := s9270;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9269; end if;
when s9270 => state := s9271; 	--9
	mulfpsclr <= '0';
when s9271 => state := s9272; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9272 => 			--11
	if (mulfprdy = '1') then state := s9273;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9272; end if;
when s9273 => state := s9274; 	--12
	mulfpsclr <= '0';
when s9274 => state := s9275; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9275 => 			--14
	if (addfprdy = '1') then state := s9276;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9275; end if;
when s9276 => state := s9277; 	--15
	addfpsclr <= '0';
when s9277 => state := s9278; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9278 => 			--17
	if (addfprdy = '1') then state := s9279;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9278; end if;
when s9279 => state := s9280; 	--18
	addfpsclr <= '0';
when s9280 => state := s9281; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9281 => 			--20
	if (addfprdy = '1') then state := s9282;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9281; end if;
when s9282 => state := s9283; 	--21
	addfpsclr <= '0';
when s9283 => state := s9284; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (477, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9284 => state := s9285; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (892, 12)); -- offset LSB 844
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s9285 => state := s9286;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (893, 12)); -- offset MSB 845
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9286 => state := s9287; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9287 => 			--4
	if (fixed2floatrdy = '1') then state := s9288;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9287; end if;
when s9288 => state := s9289; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9289 => 			--6
	if (mulfprdy = '1') then state := s9290;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9289; end if;
when s9290 => state := s9291; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9291 => 			--8
	if (mulfprdy = '1') then state := s9292;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9291; end if;
when s9292 => state := s9293; 	--9
	mulfpsclr <= '0';
when s9293 => state := s9294; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9294 => 			--11
	if (mulfprdy = '1') then state := s9295;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9294; end if;
when s9295 => state := s9296; 	--12
	mulfpsclr <= '0';
when s9296 => state := s9297; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9297 => 			--14
	if (addfprdy = '1') then state := s9298;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9297; end if;
when s9298 => state := s9299; 	--15
	addfpsclr <= '0';
when s9299 => state := s9300; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9300 => 			--17
	if (addfprdy = '1') then state := s9301;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9300; end if;
when s9301 => state := s9302; 	--18
	addfpsclr <= '0';
when s9302 => state := s9303; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9303 => 			--20
	if (addfprdy = '1') then state := s9304;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9303; end if;
when s9304 => state := s9305; 	--21
	addfpsclr <= '0';
when s9305 => state := s9306; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (478, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9306 => state := s9307; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (894, 12)); -- offset LSB 846
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s9307 => state := s9308;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (895, 12)); -- offset MSB 847
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9308 => state := s9309; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9309 => 			--4
	if (fixed2floatrdy = '1') then state := s9310;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9309; end if;
when s9310 => state := s9311; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9311 => 			--6
	if (mulfprdy = '1') then state := s9312;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9311; end if;
when s9312 => state := s9313; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9313 => 			--8
	if (mulfprdy = '1') then state := s9314;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9313; end if;
when s9314 => state := s9315; 	--9
	mulfpsclr <= '0';
when s9315 => state := s9316; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9316 => 			--11
	if (mulfprdy = '1') then state := s9317;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9316; end if;
when s9317 => state := s9318; 	--12
	mulfpsclr <= '0';
when s9318 => state := s9319; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9319 => 			--14
	if (addfprdy = '1') then state := s9320;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9319; end if;
when s9320 => state := s9321; 	--15
	addfpsclr <= '0';
when s9321 => state := s9322; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9322 => 			--17
	if (addfprdy = '1') then state := s9323;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9322; end if;
when s9323 => state := s9324; 	--18
	addfpsclr <= '0';
when s9324 => state := s9325; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9325 => 			--20
	if (addfprdy = '1') then state := s9326;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9325; end if;
when s9326 => state := s9327; 	--21
	addfpsclr <= '0';
when s9327 => state := s9328; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (479, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9328 => state := s9329; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (896, 12)); -- offset LSB 848
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s9329 => state := s9330;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (897, 12)); -- offset MSB 849
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9330 => state := s9331; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9331 => 			--4
	if (fixed2floatrdy = '1') then state := s9332;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9331; end if;
when s9332 => state := s9333; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9333 => 			--6
	if (mulfprdy = '1') then state := s9334;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9333; end if;
when s9334 => state := s9335; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9335 => 			--8
	if (mulfprdy = '1') then state := s9336;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9335; end if;
when s9336 => state := s9337; 	--9
	mulfpsclr <= '0';
when s9337 => state := s9338; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9338 => 			--11
	if (mulfprdy = '1') then state := s9339;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9338; end if;
when s9339 => state := s9340; 	--12
	mulfpsclr <= '0';
when s9340 => state := s9341; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9341 => 			--14
	if (addfprdy = '1') then state := s9342;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9341; end if;
when s9342 => state := s9343; 	--15
	addfpsclr <= '0';
when s9343 => state := s9344; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9344 => 			--17
	if (addfprdy = '1') then state := s9345;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9344; end if;
when s9345 => state := s9346; 	--18
	addfpsclr <= '0';
when s9346 => state := s9347; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9347 => 			--20
	if (addfprdy = '1') then state := s9348;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9347; end if;
when s9348 => state := s9349; 	--21
	addfpsclr <= '0';
when s9349 => state := s9350; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (480, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9350 => state := s9351; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (898, 12)); -- offset LSB 850
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s9351 => state := s9352;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (899, 12)); -- offset MSB 851
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9352 => state := s9353; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9353 => 			--4
	if (fixed2floatrdy = '1') then state := s9354;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9353; end if;
when s9354 => state := s9355; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9355 => 			--6
	if (mulfprdy = '1') then state := s9356;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9355; end if;
when s9356 => state := s9357; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9357 => 			--8
	if (mulfprdy = '1') then state := s9358;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9357; end if;
when s9358 => state := s9359; 	--9
	mulfpsclr <= '0';
when s9359 => state := s9360; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9360 => 			--11
	if (mulfprdy = '1') then state := s9361;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9360; end if;
when s9361 => state := s9362; 	--12
	mulfpsclr <= '0';
when s9362 => state := s9363; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9363 => 			--14
	if (addfprdy = '1') then state := s9364;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9363; end if;
when s9364 => state := s9365; 	--15
	addfpsclr <= '0';
when s9365 => state := s9366; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9366 => 			--17
	if (addfprdy = '1') then state := s9367;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9366; end if;
when s9367 => state := s9368; 	--18
	addfpsclr <= '0';
when s9368 => state := s9369; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9369 => 			--20
	if (addfprdy = '1') then state := s9370;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9369; end if;
when s9370 => state := s9371; 	--21
	addfpsclr <= '0';
when s9371 => state := s9372; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (481, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9372 => state := s9373; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (900, 12)); -- offset LSB 852
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s9373 => state := s9374;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (901, 12)); -- offset MSB 853
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9374 => state := s9375; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9375 => 			--4
	if (fixed2floatrdy = '1') then state := s9376;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9375; end if;
when s9376 => state := s9377; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9377 => 			--6
	if (mulfprdy = '1') then state := s9378;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9377; end if;
when s9378 => state := s9379; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9379 => 			--8
	if (mulfprdy = '1') then state := s9380;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9379; end if;
when s9380 => state := s9381; 	--9
	mulfpsclr <= '0';
when s9381 => state := s9382; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9382 => 			--11
	if (mulfprdy = '1') then state := s9383;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9382; end if;
when s9383 => state := s9384; 	--12
	mulfpsclr <= '0';
when s9384 => state := s9385; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9385 => 			--14
	if (addfprdy = '1') then state := s9386;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9385; end if;
when s9386 => state := s9387; 	--15
	addfpsclr <= '0';
when s9387 => state := s9388; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9388 => 			--17
	if (addfprdy = '1') then state := s9389;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9388; end if;
when s9389 => state := s9390; 	--18
	addfpsclr <= '0';
when s9390 => state := s9391; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9391 => 			--20
	if (addfprdy = '1') then state := s9392;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9391; end if;
when s9392 => state := s9393; 	--21
	addfpsclr <= '0';
when s9393 => state := s9394; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (482, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9394 => state := s9395; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (902, 12)); -- offset LSB 854
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s9395 => state := s9396;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (903, 12)); -- offset MSB 855
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9396 => state := s9397; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9397 => 			--4
	if (fixed2floatrdy = '1') then state := s9398;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9397; end if;
when s9398 => state := s9399; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9399 => 			--6
	if (mulfprdy = '1') then state := s9400;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9399; end if;
when s9400 => state := s9401; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9401 => 			--8
	if (mulfprdy = '1') then state := s9402;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9401; end if;
when s9402 => state := s9403; 	--9
	mulfpsclr <= '0';
when s9403 => state := s9404; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9404 => 			--11
	if (mulfprdy = '1') then state := s9405;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9404; end if;
when s9405 => state := s9406; 	--12
	mulfpsclr <= '0';
when s9406 => state := s9407; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9407 => 			--14
	if (addfprdy = '1') then state := s9408;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9407; end if;
when s9408 => state := s9409; 	--15
	addfpsclr <= '0';
when s9409 => state := s9410; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9410 => 			--17
	if (addfprdy = '1') then state := s9411;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9410; end if;
when s9411 => state := s9412; 	--18
	addfpsclr <= '0';
when s9412 => state := s9413; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9413 => 			--20
	if (addfprdy = '1') then state := s9414;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9413; end if;
when s9414 => state := s9415; 	--21
	addfpsclr <= '0';
when s9415 => state := s9416; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (483, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9416 => state := s9417; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (904, 12)); -- offset LSB 856
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s9417 => state := s9418;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (905, 12)); -- offset MSB 857
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9418 => state := s9419; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9419 => 			--4
	if (fixed2floatrdy = '1') then state := s9420;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9419; end if;
when s9420 => state := s9421; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9421 => 			--6
	if (mulfprdy = '1') then state := s9422;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9421; end if;
when s9422 => state := s9423; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9423 => 			--8
	if (mulfprdy = '1') then state := s9424;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9423; end if;
when s9424 => state := s9425; 	--9
	mulfpsclr <= '0';
when s9425 => state := s9426; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9426 => 			--11
	if (mulfprdy = '1') then state := s9427;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9426; end if;
when s9427 => state := s9428; 	--12
	mulfpsclr <= '0';
when s9428 => state := s9429; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9429 => 			--14
	if (addfprdy = '1') then state := s9430;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9429; end if;
when s9430 => state := s9431; 	--15
	addfpsclr <= '0';
when s9431 => state := s9432; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9432 => 			--17
	if (addfprdy = '1') then state := s9433;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9432; end if;
when s9433 => state := s9434; 	--18
	addfpsclr <= '0';
when s9434 => state := s9435; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9435 => 			--20
	if (addfprdy = '1') then state := s9436;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9435; end if;
when s9436 => state := s9437; 	--21
	addfpsclr <= '0';
when s9437 => state := s9438; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (484, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9438 => state := s9439; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (906, 12)); -- offset LSB 858
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s9439 => state := s9440;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (907, 12)); -- offset MSB 859
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9440 => state := s9441; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9441 => 			--4
	if (fixed2floatrdy = '1') then state := s9442;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9441; end if;
when s9442 => state := s9443; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9443 => 			--6
	if (mulfprdy = '1') then state := s9444;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9443; end if;
when s9444 => state := s9445; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9445 => 			--8
	if (mulfprdy = '1') then state := s9446;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9445; end if;
when s9446 => state := s9447; 	--9
	mulfpsclr <= '0';
when s9447 => state := s9448; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9448 => 			--11
	if (mulfprdy = '1') then state := s9449;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9448; end if;
when s9449 => state := s9450; 	--12
	mulfpsclr <= '0';
when s9450 => state := s9451; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9451 => 			--14
	if (addfprdy = '1') then state := s9452;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9451; end if;
when s9452 => state := s9453; 	--15
	addfpsclr <= '0';
when s9453 => state := s9454; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9454 => 			--17
	if (addfprdy = '1') then state := s9455;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9454; end if;
when s9455 => state := s9456; 	--18
	addfpsclr <= '0';
when s9456 => state := s9457; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9457 => 			--20
	if (addfprdy = '1') then state := s9458;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9457; end if;
when s9458 => state := s9459; 	--21
	addfpsclr <= '0';
when s9459 => state := s9460; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (485, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9460 => state := s9461; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (908, 12)); -- offset LSB 860
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s9461 => state := s9462;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (909, 12)); -- offset MSB 861
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9462 => state := s9463; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9463 => 			--4
	if (fixed2floatrdy = '1') then state := s9464;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9463; end if;
when s9464 => state := s9465; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9465 => 			--6
	if (mulfprdy = '1') then state := s9466;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9465; end if;
when s9466 => state := s9467; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9467 => 			--8
	if (mulfprdy = '1') then state := s9468;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9467; end if;
when s9468 => state := s9469; 	--9
	mulfpsclr <= '0';
when s9469 => state := s9470; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9470 => 			--11
	if (mulfprdy = '1') then state := s9471;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9470; end if;
when s9471 => state := s9472; 	--12
	mulfpsclr <= '0';
when s9472 => state := s9473; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9473 => 			--14
	if (addfprdy = '1') then state := s9474;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9473; end if;
when s9474 => state := s9475; 	--15
	addfpsclr <= '0';
when s9475 => state := s9476; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9476 => 			--17
	if (addfprdy = '1') then state := s9477;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9476; end if;
when s9477 => state := s9478; 	--18
	addfpsclr <= '0';
when s9478 => state := s9479; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9479 => 			--20
	if (addfprdy = '1') then state := s9480;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9479; end if;
when s9480 => state := s9481; 	--21
	addfpsclr <= '0';
when s9481 => state := s9482; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (486, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9482 => state := s9483; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (910, 12)); -- offset LSB 862
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s9483 => state := s9484;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (911, 12)); -- offset MSB 863
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9484 => state := s9485; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9485 => 			--4
	if (fixed2floatrdy = '1') then state := s9486;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9485; end if;
when s9486 => state := s9487; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9487 => 			--6
	if (mulfprdy = '1') then state := s9488;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9487; end if;
when s9488 => state := s9489; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9489 => 			--8
	if (mulfprdy = '1') then state := s9490;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9489; end if;
when s9490 => state := s9491; 	--9
	mulfpsclr <= '0';
when s9491 => state := s9492; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9492 => 			--11
	if (mulfprdy = '1') then state := s9493;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9492; end if;
when s9493 => state := s9494; 	--12
	mulfpsclr <= '0';
when s9494 => state := s9495; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9495 => 			--14
	if (addfprdy = '1') then state := s9496;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9495; end if;
when s9496 => state := s9497; 	--15
	addfpsclr <= '0';
when s9497 => state := s9498; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9498 => 			--17
	if (addfprdy = '1') then state := s9499;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9498; end if;
when s9499 => state := s9500; 	--18
	addfpsclr <= '0';
when s9500 => state := s9501; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9501 => 			--20
	if (addfprdy = '1') then state := s9502;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9501; end if;
when s9502 => state := s9503; 	--21
	addfpsclr <= '0';
when s9503 => state := s9504; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (487, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9504 => state := s9505; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (912, 12)); -- offset LSB 864
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s9505 => state := s9506;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (913, 12)); -- offset MSB 865
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9506 => state := s9507; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9507 => 			--4
	if (fixed2floatrdy = '1') then state := s9508;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9507; end if;
when s9508 => state := s9509; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9509 => 			--6
	if (mulfprdy = '1') then state := s9510;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9509; end if;
when s9510 => state := s9511; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9511 => 			--8
	if (mulfprdy = '1') then state := s9512;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9511; end if;
when s9512 => state := s9513; 	--9
	mulfpsclr <= '0';
when s9513 => state := s9514; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9514 => 			--11
	if (mulfprdy = '1') then state := s9515;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9514; end if;
when s9515 => state := s9516; 	--12
	mulfpsclr <= '0';
when s9516 => state := s9517; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9517 => 			--14
	if (addfprdy = '1') then state := s9518;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9517; end if;
when s9518 => state := s9519; 	--15
	addfpsclr <= '0';
when s9519 => state := s9520; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9520 => 			--17
	if (addfprdy = '1') then state := s9521;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9520; end if;
when s9521 => state := s9522; 	--18
	addfpsclr <= '0';
when s9522 => state := s9523; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9523 => 			--20
	if (addfprdy = '1') then state := s9524;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9523; end if;
when s9524 => state := s9525; 	--21
	addfpsclr <= '0';
when s9525 => state := s9526; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (488, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9526 => state := s9527; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (914, 12)); -- offset LSB 866
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s9527 => state := s9528;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (915, 12)); -- offset MSB 867
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9528 => state := s9529; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9529 => 			--4
	if (fixed2floatrdy = '1') then state := s9530;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9529; end if;
when s9530 => state := s9531; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9531 => 			--6
	if (mulfprdy = '1') then state := s9532;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9531; end if;
when s9532 => state := s9533; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9533 => 			--8
	if (mulfprdy = '1') then state := s9534;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9533; end if;
when s9534 => state := s9535; 	--9
	mulfpsclr <= '0';
when s9535 => state := s9536; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9536 => 			--11
	if (mulfprdy = '1') then state := s9537;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9536; end if;
when s9537 => state := s9538; 	--12
	mulfpsclr <= '0';
when s9538 => state := s9539; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9539 => 			--14
	if (addfprdy = '1') then state := s9540;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9539; end if;
when s9540 => state := s9541; 	--15
	addfpsclr <= '0';
when s9541 => state := s9542; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9542 => 			--17
	if (addfprdy = '1') then state := s9543;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9542; end if;
when s9543 => state := s9544; 	--18
	addfpsclr <= '0';
when s9544 => state := s9545; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9545 => 			--20
	if (addfprdy = '1') then state := s9546;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9545; end if;
when s9546 => state := s9547; 	--21
	addfpsclr <= '0';
when s9547 => state := s9548; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (489, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9548 => state := s9549; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (916, 12)); -- offset LSB 868
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s9549 => state := s9550;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (917, 12)); -- offset MSB 869
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9550 => state := s9551; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9551 => 			--4
	if (fixed2floatrdy = '1') then state := s9552;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9551; end if;
when s9552 => state := s9553; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9553 => 			--6
	if (mulfprdy = '1') then state := s9554;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9553; end if;
when s9554 => state := s9555; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9555 => 			--8
	if (mulfprdy = '1') then state := s9556;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9555; end if;
when s9556 => state := s9557; 	--9
	mulfpsclr <= '0';
when s9557 => state := s9558; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9558 => 			--11
	if (mulfprdy = '1') then state := s9559;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9558; end if;
when s9559 => state := s9560; 	--12
	mulfpsclr <= '0';
when s9560 => state := s9561; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9561 => 			--14
	if (addfprdy = '1') then state := s9562;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9561; end if;
when s9562 => state := s9563; 	--15
	addfpsclr <= '0';
when s9563 => state := s9564; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9564 => 			--17
	if (addfprdy = '1') then state := s9565;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9564; end if;
when s9565 => state := s9566; 	--18
	addfpsclr <= '0';
when s9566 => state := s9567; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9567 => 			--20
	if (addfprdy = '1') then state := s9568;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9567; end if;
when s9568 => state := s9569; 	--21
	addfpsclr <= '0';
when s9569 => state := s9570; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (490, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9570 => state := s9571; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (918, 12)); -- offset LSB 870
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s9571 => state := s9572;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (919, 12)); -- offset MSB 871
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9572 => state := s9573; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9573 => 			--4
	if (fixed2floatrdy = '1') then state := s9574;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9573; end if;
when s9574 => state := s9575; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9575 => 			--6
	if (mulfprdy = '1') then state := s9576;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9575; end if;
when s9576 => state := s9577; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9577 => 			--8
	if (mulfprdy = '1') then state := s9578;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9577; end if;
when s9578 => state := s9579; 	--9
	mulfpsclr <= '0';
when s9579 => state := s9580; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9580 => 			--11
	if (mulfprdy = '1') then state := s9581;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9580; end if;
when s9581 => state := s9582; 	--12
	mulfpsclr <= '0';
when s9582 => state := s9583; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9583 => 			--14
	if (addfprdy = '1') then state := s9584;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9583; end if;
when s9584 => state := s9585; 	--15
	addfpsclr <= '0';
when s9585 => state := s9586; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9586 => 			--17
	if (addfprdy = '1') then state := s9587;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9586; end if;
when s9587 => state := s9588; 	--18
	addfpsclr <= '0';
when s9588 => state := s9589; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9589 => 			--20
	if (addfprdy = '1') then state := s9590;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9589; end if;
when s9590 => state := s9591; 	--21
	addfpsclr <= '0';
when s9591 => state := s9592; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (491, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9592 => state := s9593; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (920, 12)); -- offset LSB 872
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s9593 => state := s9594;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (921, 12)); -- offset MSB 873
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9594 => state := s9595; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9595 => 			--4
	if (fixed2floatrdy = '1') then state := s9596;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9595; end if;
when s9596 => state := s9597; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9597 => 			--6
	if (mulfprdy = '1') then state := s9598;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9597; end if;
when s9598 => state := s9599; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9599 => 			--8
	if (mulfprdy = '1') then state := s9600;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9599; end if;
when s9600 => state := s9601; 	--9
	mulfpsclr <= '0';
when s9601 => state := s9602; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9602 => 			--11
	if (mulfprdy = '1') then state := s9603;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9602; end if;
when s9603 => state := s9604; 	--12
	mulfpsclr <= '0';
when s9604 => state := s9605; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9605 => 			--14
	if (addfprdy = '1') then state := s9606;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9605; end if;
when s9606 => state := s9607; 	--15
	addfpsclr <= '0';
when s9607 => state := s9608; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9608 => 			--17
	if (addfprdy = '1') then state := s9609;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9608; end if;
when s9609 => state := s9610; 	--18
	addfpsclr <= '0';
when s9610 => state := s9611; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9611 => 			--20
	if (addfprdy = '1') then state := s9612;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9611; end if;
when s9612 => state := s9613; 	--21
	addfpsclr <= '0';
when s9613 => state := s9614; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (492, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9614 => state := s9615; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (922, 12)); -- offset LSB 874
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s9615 => state := s9616;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (923, 12)); -- offset MSB 875
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9616 => state := s9617; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9617 => 			--4
	if (fixed2floatrdy = '1') then state := s9618;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9617; end if;
when s9618 => state := s9619; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9619 => 			--6
	if (mulfprdy = '1') then state := s9620;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9619; end if;
when s9620 => state := s9621; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9621 => 			--8
	if (mulfprdy = '1') then state := s9622;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9621; end if;
when s9622 => state := s9623; 	--9
	mulfpsclr <= '0';
when s9623 => state := s9624; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9624 => 			--11
	if (mulfprdy = '1') then state := s9625;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9624; end if;
when s9625 => state := s9626; 	--12
	mulfpsclr <= '0';
when s9626 => state := s9627; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9627 => 			--14
	if (addfprdy = '1') then state := s9628;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9627; end if;
when s9628 => state := s9629; 	--15
	addfpsclr <= '0';
when s9629 => state := s9630; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9630 => 			--17
	if (addfprdy = '1') then state := s9631;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9630; end if;
when s9631 => state := s9632; 	--18
	addfpsclr <= '0';
when s9632 => state := s9633; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9633 => 			--20
	if (addfprdy = '1') then state := s9634;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9633; end if;
when s9634 => state := s9635; 	--21
	addfpsclr <= '0';
when s9635 => state := s9636; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (493, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9636 => state := s9637; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (924, 12)); -- offset LSB 876
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s9637 => state := s9638;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (925, 12)); -- offset MSB 877
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9638 => state := s9639; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9639 => 			--4
	if (fixed2floatrdy = '1') then state := s9640;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9639; end if;
when s9640 => state := s9641; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9641 => 			--6
	if (mulfprdy = '1') then state := s9642;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9641; end if;
when s9642 => state := s9643; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9643 => 			--8
	if (mulfprdy = '1') then state := s9644;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9643; end if;
when s9644 => state := s9645; 	--9
	mulfpsclr <= '0';
when s9645 => state := s9646; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9646 => 			--11
	if (mulfprdy = '1') then state := s9647;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9646; end if;
when s9647 => state := s9648; 	--12
	mulfpsclr <= '0';
when s9648 => state := s9649; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9649 => 			--14
	if (addfprdy = '1') then state := s9650;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9649; end if;
when s9650 => state := s9651; 	--15
	addfpsclr <= '0';
when s9651 => state := s9652; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9652 => 			--17
	if (addfprdy = '1') then state := s9653;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9652; end if;
when s9653 => state := s9654; 	--18
	addfpsclr <= '0';
when s9654 => state := s9655; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9655 => 			--20
	if (addfprdy = '1') then state := s9656;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9655; end if;
when s9656 => state := s9657; 	--21
	addfpsclr <= '0';
when s9657 => state := s9658; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (494, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9658 => state := s9659; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (926, 12)); -- offset LSB 878
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s9659 => state := s9660;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (927, 12)); -- offset MSB 879
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9660 => state := s9661; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9661 => 			--4
	if (fixed2floatrdy = '1') then state := s9662;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9661; end if;
when s9662 => state := s9663; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9663 => 			--6
	if (mulfprdy = '1') then state := s9664;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9663; end if;
when s9664 => state := s9665; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9665 => 			--8
	if (mulfprdy = '1') then state := s9666;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9665; end if;
when s9666 => state := s9667; 	--9
	mulfpsclr <= '0';
when s9667 => state := s9668; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9668 => 			--11
	if (mulfprdy = '1') then state := s9669;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9668; end if;
when s9669 => state := s9670; 	--12
	mulfpsclr <= '0';
when s9670 => state := s9671; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9671 => 			--14
	if (addfprdy = '1') then state := s9672;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9671; end if;
when s9672 => state := s9673; 	--15
	addfpsclr <= '0';
when s9673 => state := s9674; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9674 => 			--17
	if (addfprdy = '1') then state := s9675;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9674; end if;
when s9675 => state := s9676; 	--18
	addfpsclr <= '0';
when s9676 => state := s9677; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9677 => 			--20
	if (addfprdy = '1') then state := s9678;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9677; end if;
when s9678 => state := s9679; 	--21
	addfpsclr <= '0';
when s9679 => state := s9680; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (495, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9680 => state := s9681; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (928, 12)); -- offset LSB 880
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s9681 => state := s9682;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (929, 12)); -- offset MSB 881
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9682 => state := s9683; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9683 => 			--4
	if (fixed2floatrdy = '1') then state := s9684;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9683; end if;
when s9684 => state := s9685; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9685 => 			--6
	if (mulfprdy = '1') then state := s9686;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9685; end if;
when s9686 => state := s9687; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9687 => 			--8
	if (mulfprdy = '1') then state := s9688;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9687; end if;
when s9688 => state := s9689; 	--9
	mulfpsclr <= '0';
when s9689 => state := s9690; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9690 => 			--11
	if (mulfprdy = '1') then state := s9691;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9690; end if;
when s9691 => state := s9692; 	--12
	mulfpsclr <= '0';
when s9692 => state := s9693; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9693 => 			--14
	if (addfprdy = '1') then state := s9694;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9693; end if;
when s9694 => state := s9695; 	--15
	addfpsclr <= '0';
when s9695 => state := s9696; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9696 => 			--17
	if (addfprdy = '1') then state := s9697;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9696; end if;
when s9697 => state := s9698; 	--18
	addfpsclr <= '0';
when s9698 => state := s9699; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9699 => 			--20
	if (addfprdy = '1') then state := s9700;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9699; end if;
when s9700 => state := s9701; 	--21
	addfpsclr <= '0';
when s9701 => state := s9702; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (496, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9702 => state := s9703; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (930, 12)); -- offset LSB 882
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s9703 => state := s9704;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (931, 12)); -- offset MSB 883
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9704 => state := s9705; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9705 => 			--4
	if (fixed2floatrdy = '1') then state := s9706;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9705; end if;
when s9706 => state := s9707; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9707 => 			--6
	if (mulfprdy = '1') then state := s9708;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9707; end if;
when s9708 => state := s9709; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9709 => 			--8
	if (mulfprdy = '1') then state := s9710;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9709; end if;
when s9710 => state := s9711; 	--9
	mulfpsclr <= '0';
when s9711 => state := s9712; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9712 => 			--11
	if (mulfprdy = '1') then state := s9713;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9712; end if;
when s9713 => state := s9714; 	--12
	mulfpsclr <= '0';
when s9714 => state := s9715; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9715 => 			--14
	if (addfprdy = '1') then state := s9716;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9715; end if;
when s9716 => state := s9717; 	--15
	addfpsclr <= '0';
when s9717 => state := s9718; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9718 => 			--17
	if (addfprdy = '1') then state := s9719;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9718; end if;
when s9719 => state := s9720; 	--18
	addfpsclr <= '0';
when s9720 => state := s9721; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9721 => 			--20
	if (addfprdy = '1') then state := s9722;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9721; end if;
when s9722 => state := s9723; 	--21
	addfpsclr <= '0';
when s9723 => state := s9724; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (497, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9724 => state := s9725; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (932, 12)); -- offset LSB 884
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s9725 => state := s9726;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (933, 12)); -- offset MSB 885
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9726 => state := s9727; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9727 => 			--4
	if (fixed2floatrdy = '1') then state := s9728;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9727; end if;
when s9728 => state := s9729; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9729 => 			--6
	if (mulfprdy = '1') then state := s9730;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9729; end if;
when s9730 => state := s9731; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9731 => 			--8
	if (mulfprdy = '1') then state := s9732;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9731; end if;
when s9732 => state := s9733; 	--9
	mulfpsclr <= '0';
when s9733 => state := s9734; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9734 => 			--11
	if (mulfprdy = '1') then state := s9735;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9734; end if;
when s9735 => state := s9736; 	--12
	mulfpsclr <= '0';
when s9736 => state := s9737; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9737 => 			--14
	if (addfprdy = '1') then state := s9738;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9737; end if;
when s9738 => state := s9739; 	--15
	addfpsclr <= '0';
when s9739 => state := s9740; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9740 => 			--17
	if (addfprdy = '1') then state := s9741;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9740; end if;
when s9741 => state := s9742; 	--18
	addfpsclr <= '0';
when s9742 => state := s9743; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9743 => 			--20
	if (addfprdy = '1') then state := s9744;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9743; end if;
when s9744 => state := s9745; 	--21
	addfpsclr <= '0';
when s9745 => state := s9746; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (498, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9746 => state := s9747; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (934, 12)); -- offset LSB 886
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s9747 => state := s9748;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (935, 12)); -- offset MSB 887
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9748 => state := s9749; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9749 => 			--4
	if (fixed2floatrdy = '1') then state := s9750;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9749; end if;
when s9750 => state := s9751; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9751 => 			--6
	if (mulfprdy = '1') then state := s9752;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9751; end if;
when s9752 => state := s9753; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9753 => 			--8
	if (mulfprdy = '1') then state := s9754;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9753; end if;
when s9754 => state := s9755; 	--9
	mulfpsclr <= '0';
when s9755 => state := s9756; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9756 => 			--11
	if (mulfprdy = '1') then state := s9757;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9756; end if;
when s9757 => state := s9758; 	--12
	mulfpsclr <= '0';
when s9758 => state := s9759; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9759 => 			--14
	if (addfprdy = '1') then state := s9760;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9759; end if;
when s9760 => state := s9761; 	--15
	addfpsclr <= '0';
when s9761 => state := s9762; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9762 => 			--17
	if (addfprdy = '1') then state := s9763;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9762; end if;
when s9763 => state := s9764; 	--18
	addfpsclr <= '0';
when s9764 => state := s9765; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9765 => 			--20
	if (addfprdy = '1') then state := s9766;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9765; end if;
when s9766 => state := s9767; 	--21
	addfpsclr <= '0';
when s9767 => state := s9768; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (499, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9768 => state := s9769; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (936, 12)); -- offset LSB 888
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s9769 => state := s9770;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (937, 12)); -- offset MSB 889
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9770 => state := s9771; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9771 => 			--4
	if (fixed2floatrdy = '1') then state := s9772;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9771; end if;
when s9772 => state := s9773; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9773 => 			--6
	if (mulfprdy = '1') then state := s9774;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9773; end if;
when s9774 => state := s9775; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9775 => 			--8
	if (mulfprdy = '1') then state := s9776;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9775; end if;
when s9776 => state := s9777; 	--9
	mulfpsclr <= '0';
when s9777 => state := s9778; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9778 => 			--11
	if (mulfprdy = '1') then state := s9779;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9778; end if;
when s9779 => state := s9780; 	--12
	mulfpsclr <= '0';
when s9780 => state := s9781; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9781 => 			--14
	if (addfprdy = '1') then state := s9782;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9781; end if;
when s9782 => state := s9783; 	--15
	addfpsclr <= '0';
when s9783 => state := s9784; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9784 => 			--17
	if (addfprdy = '1') then state := s9785;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9784; end if;
when s9785 => state := s9786; 	--18
	addfpsclr <= '0';
when s9786 => state := s9787; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9787 => 			--20
	if (addfprdy = '1') then state := s9788;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9787; end if;
when s9788 => state := s9789; 	--21
	addfpsclr <= '0';
when s9789 => state := s9790; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (500, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9790 => state := s9791; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (938, 12)); -- offset LSB 890
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s9791 => state := s9792;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (939, 12)); -- offset MSB 891
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9792 => state := s9793; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9793 => 			--4
	if (fixed2floatrdy = '1') then state := s9794;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9793; end if;
when s9794 => state := s9795; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9795 => 			--6
	if (mulfprdy = '1') then state := s9796;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9795; end if;
when s9796 => state := s9797; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9797 => 			--8
	if (mulfprdy = '1') then state := s9798;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9797; end if;
when s9798 => state := s9799; 	--9
	mulfpsclr <= '0';
when s9799 => state := s9800; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9800 => 			--11
	if (mulfprdy = '1') then state := s9801;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9800; end if;
when s9801 => state := s9802; 	--12
	mulfpsclr <= '0';
when s9802 => state := s9803; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9803 => 			--14
	if (addfprdy = '1') then state := s9804;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9803; end if;
when s9804 => state := s9805; 	--15
	addfpsclr <= '0';
when s9805 => state := s9806; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9806 => 			--17
	if (addfprdy = '1') then state := s9807;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9806; end if;
when s9807 => state := s9808; 	--18
	addfpsclr <= '0';
when s9808 => state := s9809; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9809 => 			--20
	if (addfprdy = '1') then state := s9810;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9809; end if;
when s9810 => state := s9811; 	--21
	addfpsclr <= '0';
when s9811 => state := s9812; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (501, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9812 => state := s9813; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (940, 12)); -- offset LSB 892
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s9813 => state := s9814;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (941, 12)); -- offset MSB 893
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9814 => state := s9815; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9815 => 			--4
	if (fixed2floatrdy = '1') then state := s9816;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9815; end if;
when s9816 => state := s9817; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9817 => 			--6
	if (mulfprdy = '1') then state := s9818;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9817; end if;
when s9818 => state := s9819; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9819 => 			--8
	if (mulfprdy = '1') then state := s9820;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9819; end if;
when s9820 => state := s9821; 	--9
	mulfpsclr <= '0';
when s9821 => state := s9822; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9822 => 			--11
	if (mulfprdy = '1') then state := s9823;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9822; end if;
when s9823 => state := s9824; 	--12
	mulfpsclr <= '0';
when s9824 => state := s9825; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9825 => 			--14
	if (addfprdy = '1') then state := s9826;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9825; end if;
when s9826 => state := s9827; 	--15
	addfpsclr <= '0';
when s9827 => state := s9828; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9828 => 			--17
	if (addfprdy = '1') then state := s9829;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9828; end if;
when s9829 => state := s9830; 	--18
	addfpsclr <= '0';
when s9830 => state := s9831; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9831 => 			--20
	if (addfprdy = '1') then state := s9832;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9831; end if;
when s9832 => state := s9833; 	--21
	addfpsclr <= '0';
when s9833 => state := s9834; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (502, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9834 => state := s9835; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (942, 12)); -- offset LSB 894
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s9835 => state := s9836;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (943, 12)); -- offset MSB 895
	addra <= std_logic_vector (to_unsigned (13, 10)); -- OCCrowI 13
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9836 => state := s9837; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9837 => 			--4
	if (fixed2floatrdy = '1') then state := s9838;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9837; end if;
when s9838 => state := s9839; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9839 => 			--6
	if (mulfprdy = '1') then state := s9840;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9839; end if;
when s9840 => state := s9841; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9841 => 			--8
	if (mulfprdy = '1') then state := s9842;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9841; end if;
when s9842 => state := s9843; 	--9
	mulfpsclr <= '0';
when s9843 => state := s9844; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9844 => 			--11
	if (mulfprdy = '1') then state := s9845;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9844; end if;
when s9845 => state := s9846; 	--12
	mulfpsclr <= '0';
when s9846 => state := s9847; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9847 => 			--14
	if (addfprdy = '1') then state := s9848;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9847; end if;
when s9848 => state := s9849; 	--15
	addfpsclr <= '0';
when s9849 => state := s9850; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9850 => 			--17
	if (addfprdy = '1') then state := s9851;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9850; end if;
when s9851 => state := s9852; 	--18
	addfpsclr <= '0';
when s9852 => state := s9853; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9853 => 			--20
	if (addfprdy = '1') then state := s9854;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9853; end if;
when s9854 => state := s9855; 	--21
	addfpsclr <= '0';
when s9855 => state := s9856; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (503, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9856 => state := s9857; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (944, 12)); -- offset LSB 896
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s9857 => state := s9858;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (945, 12)); -- offset MSB 897
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9858 => state := s9859; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9859 => 			--4
	if (fixed2floatrdy = '1') then state := s9860;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9859; end if;
when s9860 => state := s9861; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9861 => 			--6
	if (mulfprdy = '1') then state := s9862;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9861; end if;
when s9862 => state := s9863; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9863 => 			--8
	if (mulfprdy = '1') then state := s9864;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9863; end if;
when s9864 => state := s9865; 	--9
	mulfpsclr <= '0';
when s9865 => state := s9866; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9866 => 			--11
	if (mulfprdy = '1') then state := s9867;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9866; end if;
when s9867 => state := s9868; 	--12
	mulfpsclr <= '0';
when s9868 => state := s9869; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9869 => 			--14
	if (addfprdy = '1') then state := s9870;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9869; end if;
when s9870 => state := s9871; 	--15
	addfpsclr <= '0';
when s9871 => state := s9872; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9872 => 			--17
	if (addfprdy = '1') then state := s9873;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9872; end if;
when s9873 => state := s9874; 	--18
	addfpsclr <= '0';
when s9874 => state := s9875; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9875 => 			--20
	if (addfprdy = '1') then state := s9876;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9875; end if;
when s9876 => state := s9877; 	--21
	addfpsclr <= '0';
when s9877 => state := s9878; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (504, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9878 => state := s9879; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (946, 12)); -- offset LSB 898
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s9879 => state := s9880;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (947, 12)); -- offset MSB 899
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9880 => state := s9881; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9881 => 			--4
	if (fixed2floatrdy = '1') then state := s9882;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9881; end if;
when s9882 => state := s9883; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9883 => 			--6
	if (mulfprdy = '1') then state := s9884;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9883; end if;
when s9884 => state := s9885; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9885 => 			--8
	if (mulfprdy = '1') then state := s9886;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9885; end if;
when s9886 => state := s9887; 	--9
	mulfpsclr <= '0';
when s9887 => state := s9888; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9888 => 			--11
	if (mulfprdy = '1') then state := s9889;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9888; end if;
when s9889 => state := s9890; 	--12
	mulfpsclr <= '0';
when s9890 => state := s9891; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9891 => 			--14
	if (addfprdy = '1') then state := s9892;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9891; end if;
when s9892 => state := s9893; 	--15
	addfpsclr <= '0';
when s9893 => state := s9894; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9894 => 			--17
	if (addfprdy = '1') then state := s9895;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9894; end if;
when s9895 => state := s9896; 	--18
	addfpsclr <= '0';
when s9896 => state := s9897; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9897 => 			--20
	if (addfprdy = '1') then state := s9898;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9897; end if;
when s9898 => state := s9899; 	--21
	addfpsclr <= '0';
when s9899 => state := s9900; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (505, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9900 => state := s9901; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (948, 12)); -- offset LSB 900
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s9901 => state := s9902;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (949, 12)); -- offset MSB 901
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9902 => state := s9903; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9903 => 			--4
	if (fixed2floatrdy = '1') then state := s9904;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9903; end if;
when s9904 => state := s9905; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9905 => 			--6
	if (mulfprdy = '1') then state := s9906;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9905; end if;
when s9906 => state := s9907; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9907 => 			--8
	if (mulfprdy = '1') then state := s9908;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9907; end if;
when s9908 => state := s9909; 	--9
	mulfpsclr <= '0';
when s9909 => state := s9910; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9910 => 			--11
	if (mulfprdy = '1') then state := s9911;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9910; end if;
when s9911 => state := s9912; 	--12
	mulfpsclr <= '0';
when s9912 => state := s9913; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9913 => 			--14
	if (addfprdy = '1') then state := s9914;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9913; end if;
when s9914 => state := s9915; 	--15
	addfpsclr <= '0';
when s9915 => state := s9916; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9916 => 			--17
	if (addfprdy = '1') then state := s9917;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9916; end if;
when s9917 => state := s9918; 	--18
	addfpsclr <= '0';
when s9918 => state := s9919; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9919 => 			--20
	if (addfprdy = '1') then state := s9920;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9919; end if;
when s9920 => state := s9921; 	--21
	addfpsclr <= '0';
when s9921 => state := s9922; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (506, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9922 => state := s9923; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (950, 12)); -- offset LSB 902
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s9923 => state := s9924;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (951, 12)); -- offset MSB 903
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9924 => state := s9925; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9925 => 			--4
	if (fixed2floatrdy = '1') then state := s9926;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9925; end if;
when s9926 => state := s9927; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9927 => 			--6
	if (mulfprdy = '1') then state := s9928;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9927; end if;
when s9928 => state := s9929; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9929 => 			--8
	if (mulfprdy = '1') then state := s9930;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9929; end if;
when s9930 => state := s9931; 	--9
	mulfpsclr <= '0';
when s9931 => state := s9932; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9932 => 			--11
	if (mulfprdy = '1') then state := s9933;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9932; end if;
when s9933 => state := s9934; 	--12
	mulfpsclr <= '0';
when s9934 => state := s9935; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9935 => 			--14
	if (addfprdy = '1') then state := s9936;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9935; end if;
when s9936 => state := s9937; 	--15
	addfpsclr <= '0';
when s9937 => state := s9938; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9938 => 			--17
	if (addfprdy = '1') then state := s9939;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9938; end if;
when s9939 => state := s9940; 	--18
	addfpsclr <= '0';
when s9940 => state := s9941; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9941 => 			--20
	if (addfprdy = '1') then state := s9942;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9941; end if;
when s9942 => state := s9943; 	--21
	addfpsclr <= '0';
when s9943 => state := s9944; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (507, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9944 => state := s9945; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (952, 12)); -- offset LSB 904
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s9945 => state := s9946;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (953, 12)); -- offset MSB 905
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9946 => state := s9947; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9947 => 			--4
	if (fixed2floatrdy = '1') then state := s9948;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9947; end if;
when s9948 => state := s9949; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9949 => 			--6
	if (mulfprdy = '1') then state := s9950;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9949; end if;
when s9950 => state := s9951; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9951 => 			--8
	if (mulfprdy = '1') then state := s9952;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9951; end if;
when s9952 => state := s9953; 	--9
	mulfpsclr <= '0';
when s9953 => state := s9954; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9954 => 			--11
	if (mulfprdy = '1') then state := s9955;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9954; end if;
when s9955 => state := s9956; 	--12
	mulfpsclr <= '0';
when s9956 => state := s9957; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9957 => 			--14
	if (addfprdy = '1') then state := s9958;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9957; end if;
when s9958 => state := s9959; 	--15
	addfpsclr <= '0';
when s9959 => state := s9960; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9960 => 			--17
	if (addfprdy = '1') then state := s9961;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9960; end if;
when s9961 => state := s9962; 	--18
	addfpsclr <= '0';
when s9962 => state := s9963; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9963 => 			--20
	if (addfprdy = '1') then state := s9964;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9963; end if;
when s9964 => state := s9965; 	--21
	addfpsclr <= '0';
when s9965 => state := s9966; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (508, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9966 => state := s9967; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (954, 12)); -- offset LSB 906
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s9967 => state := s9968;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (955, 12)); -- offset MSB 907
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9968 => state := s9969; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9969 => 			--4
	if (fixed2floatrdy = '1') then state := s9970;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9969; end if;
when s9970 => state := s9971; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9971 => 			--6
	if (mulfprdy = '1') then state := s9972;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9971; end if;
when s9972 => state := s9973; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9973 => 			--8
	if (mulfprdy = '1') then state := s9974;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9973; end if;
when s9974 => state := s9975; 	--9
	mulfpsclr <= '0';
when s9975 => state := s9976; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9976 => 			--11
	if (mulfprdy = '1') then state := s9977;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9976; end if;
when s9977 => state := s9978; 	--12
	mulfpsclr <= '0';
when s9978 => state := s9979; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s9979 => 			--14
	if (addfprdy = '1') then state := s9980;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9979; end if;
when s9980 => state := s9981; 	--15
	addfpsclr <= '0';
when s9981 => state := s9982; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s9982 => 			--17
	if (addfprdy = '1') then state := s9983;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9982; end if;
when s9983 => state := s9984; 	--18
	addfpsclr <= '0';
when s9984 => state := s9985; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s9985 => 			--20
	if (addfprdy = '1') then state := s9986;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s9985; end if;
when s9986 => state := s9987; 	--21
	addfpsclr <= '0';
when s9987 => state := s9988; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (509, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s9988 => state := s9989; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (956, 12)); -- offset LSB 908
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s9989 => state := s9990;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (957, 12)); -- offset MSB 909
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s9990 => state := s9991; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s9991 => 			--4
	if (fixed2floatrdy = '1') then state := s9992;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s9991; end if;
when s9992 => state := s9993; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s9993 => 			--6
	if (mulfprdy = '1') then state := s9994;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9993; end if;
when s9994 => state := s9995; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s9995 => 			--8
	if (mulfprdy = '1') then state := s9996;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9995; end if;
when s9996 => state := s9997; 	--9
	mulfpsclr <= '0';
when s9997 => state := s9998; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s9998 => 			--11
	if (mulfprdy = '1') then state := s9999;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s9998; end if;
when s9999 => state := s10000; 	--12
	mulfpsclr <= '0';
when s10000 => state := s10001; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10001 => 			--14
	if (addfprdy = '1') then state := s10002;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10001; end if;
when s10002 => state := s10003; 	--15
	addfpsclr <= '0';
when s10003 => state := s10004; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10004 => 			--17
	if (addfprdy = '1') then state := s10005;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10004; end if;
when s10005 => state := s10006; 	--18
	addfpsclr <= '0';
when s10006 => state := s10007; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10007 => 			--20
	if (addfprdy = '1') then state := s10008;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10007; end if;
when s10008 => state := s10009; 	--21
	addfpsclr <= '0';
when s10009 => state := s10010; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (510, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10010 => state := s10011; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (958, 12)); -- offset LSB 910
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s10011 => state := s10012;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (959, 12)); -- offset MSB 911
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10012 => state := s10013; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10013 => 			--4
	if (fixed2floatrdy = '1') then state := s10014;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10013; end if;
when s10014 => state := s10015; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10015 => 			--6
	if (mulfprdy = '1') then state := s10016;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10015; end if;
when s10016 => state := s10017; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10017 => 			--8
	if (mulfprdy = '1') then state := s10018;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10017; end if;
when s10018 => state := s10019; 	--9
	mulfpsclr <= '0';
when s10019 => state := s10020; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10020 => 			--11
	if (mulfprdy = '1') then state := s10021;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10020; end if;
when s10021 => state := s10022; 	--12
	mulfpsclr <= '0';
when s10022 => state := s10023; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10023 => 			--14
	if (addfprdy = '1') then state := s10024;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10023; end if;
when s10024 => state := s10025; 	--15
	addfpsclr <= '0';
when s10025 => state := s10026; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10026 => 			--17
	if (addfprdy = '1') then state := s10027;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10026; end if;
when s10027 => state := s10028; 	--18
	addfpsclr <= '0';
when s10028 => state := s10029; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10029 => 			--20
	if (addfprdy = '1') then state := s10030;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10029; end if;
when s10030 => state := s10031; 	--21
	addfpsclr <= '0';
when s10031 => state := s10032; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (511, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10032 => state := s10033; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (960, 12)); -- offset LSB 912
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s10033 => state := s10034;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (961, 12)); -- offset MSB 913
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10034 => state := s10035; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10035 => 			--4
	if (fixed2floatrdy = '1') then state := s10036;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10035; end if;
when s10036 => state := s10037; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10037 => 			--6
	if (mulfprdy = '1') then state := s10038;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10037; end if;
when s10038 => state := s10039; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10039 => 			--8
	if (mulfprdy = '1') then state := s10040;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10039; end if;
when s10040 => state := s10041; 	--9
	mulfpsclr <= '0';
when s10041 => state := s10042; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10042 => 			--11
	if (mulfprdy = '1') then state := s10043;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10042; end if;
when s10043 => state := s10044; 	--12
	mulfpsclr <= '0';
when s10044 => state := s10045; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10045 => 			--14
	if (addfprdy = '1') then state := s10046;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10045; end if;
when s10046 => state := s10047; 	--15
	addfpsclr <= '0';
when s10047 => state := s10048; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10048 => 			--17
	if (addfprdy = '1') then state := s10049;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10048; end if;
when s10049 => state := s10050; 	--18
	addfpsclr <= '0';
when s10050 => state := s10051; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10051 => 			--20
	if (addfprdy = '1') then state := s10052;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10051; end if;
when s10052 => state := s10053; 	--21
	addfpsclr <= '0';
when s10053 => state := s10054; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (512, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10054 => state := s10055; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (962, 12)); -- offset LSB 914
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s10055 => state := s10056;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (963, 12)); -- offset MSB 915
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10056 => state := s10057; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10057 => 			--4
	if (fixed2floatrdy = '1') then state := s10058;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10057; end if;
when s10058 => state := s10059; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10059 => 			--6
	if (mulfprdy = '1') then state := s10060;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10059; end if;
when s10060 => state := s10061; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10061 => 			--8
	if (mulfprdy = '1') then state := s10062;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10061; end if;
when s10062 => state := s10063; 	--9
	mulfpsclr <= '0';
when s10063 => state := s10064; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10064 => 			--11
	if (mulfprdy = '1') then state := s10065;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10064; end if;
when s10065 => state := s10066; 	--12
	mulfpsclr <= '0';
when s10066 => state := s10067; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10067 => 			--14
	if (addfprdy = '1') then state := s10068;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10067; end if;
when s10068 => state := s10069; 	--15
	addfpsclr <= '0';
when s10069 => state := s10070; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10070 => 			--17
	if (addfprdy = '1') then state := s10071;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10070; end if;
when s10071 => state := s10072; 	--18
	addfpsclr <= '0';
when s10072 => state := s10073; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10073 => 			--20
	if (addfprdy = '1') then state := s10074;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10073; end if;
when s10074 => state := s10075; 	--21
	addfpsclr <= '0';
when s10075 => state := s10076; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (513, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10076 => state := s10077; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (964, 12)); -- offset LSB 916
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s10077 => state := s10078;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (965, 12)); -- offset MSB 917
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10078 => state := s10079; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10079 => 			--4
	if (fixed2floatrdy = '1') then state := s10080;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10079; end if;
when s10080 => state := s10081; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10081 => 			--6
	if (mulfprdy = '1') then state := s10082;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10081; end if;
when s10082 => state := s10083; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10083 => 			--8
	if (mulfprdy = '1') then state := s10084;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10083; end if;
when s10084 => state := s10085; 	--9
	mulfpsclr <= '0';
when s10085 => state := s10086; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10086 => 			--11
	if (mulfprdy = '1') then state := s10087;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10086; end if;
when s10087 => state := s10088; 	--12
	mulfpsclr <= '0';
when s10088 => state := s10089; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10089 => 			--14
	if (addfprdy = '1') then state := s10090;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10089; end if;
when s10090 => state := s10091; 	--15
	addfpsclr <= '0';
when s10091 => state := s10092; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10092 => 			--17
	if (addfprdy = '1') then state := s10093;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10092; end if;
when s10093 => state := s10094; 	--18
	addfpsclr <= '0';
when s10094 => state := s10095; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10095 => 			--20
	if (addfprdy = '1') then state := s10096;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10095; end if;
when s10096 => state := s10097; 	--21
	addfpsclr <= '0';
when s10097 => state := s10098; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (514, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10098 => state := s10099; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (966, 12)); -- offset LSB 918
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s10099 => state := s10100;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (967, 12)); -- offset MSB 919
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10100 => state := s10101; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10101 => 			--4
	if (fixed2floatrdy = '1') then state := s10102;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10101; end if;
when s10102 => state := s10103; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10103 => 			--6
	if (mulfprdy = '1') then state := s10104;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10103; end if;
when s10104 => state := s10105; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10105 => 			--8
	if (mulfprdy = '1') then state := s10106;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10105; end if;
when s10106 => state := s10107; 	--9
	mulfpsclr <= '0';
when s10107 => state := s10108; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10108 => 			--11
	if (mulfprdy = '1') then state := s10109;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10108; end if;
when s10109 => state := s10110; 	--12
	mulfpsclr <= '0';
when s10110 => state := s10111; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10111 => 			--14
	if (addfprdy = '1') then state := s10112;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10111; end if;
when s10112 => state := s10113; 	--15
	addfpsclr <= '0';
when s10113 => state := s10114; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10114 => 			--17
	if (addfprdy = '1') then state := s10115;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10114; end if;
when s10115 => state := s10116; 	--18
	addfpsclr <= '0';
when s10116 => state := s10117; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10117 => 			--20
	if (addfprdy = '1') then state := s10118;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10117; end if;
when s10118 => state := s10119; 	--21
	addfpsclr <= '0';
when s10119 => state := s10120; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (515, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10120 => state := s10121; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (968, 12)); -- offset LSB 920
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s10121 => state := s10122;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (969, 12)); -- offset MSB 921
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10122 => state := s10123; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10123 => 			--4
	if (fixed2floatrdy = '1') then state := s10124;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10123; end if;
when s10124 => state := s10125; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10125 => 			--6
	if (mulfprdy = '1') then state := s10126;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10125; end if;
when s10126 => state := s10127; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10127 => 			--8
	if (mulfprdy = '1') then state := s10128;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10127; end if;
when s10128 => state := s10129; 	--9
	mulfpsclr <= '0';
when s10129 => state := s10130; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10130 => 			--11
	if (mulfprdy = '1') then state := s10131;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10130; end if;
when s10131 => state := s10132; 	--12
	mulfpsclr <= '0';
when s10132 => state := s10133; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10133 => 			--14
	if (addfprdy = '1') then state := s10134;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10133; end if;
when s10134 => state := s10135; 	--15
	addfpsclr <= '0';
when s10135 => state := s10136; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10136 => 			--17
	if (addfprdy = '1') then state := s10137;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10136; end if;
when s10137 => state := s10138; 	--18
	addfpsclr <= '0';
when s10138 => state := s10139; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10139 => 			--20
	if (addfprdy = '1') then state := s10140;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10139; end if;
when s10140 => state := s10141; 	--21
	addfpsclr <= '0';
when s10141 => state := s10142; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (516, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10142 => state := s10143; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (970, 12)); -- offset LSB 922
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s10143 => state := s10144;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (971, 12)); -- offset MSB 923
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10144 => state := s10145; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10145 => 			--4
	if (fixed2floatrdy = '1') then state := s10146;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10145; end if;
when s10146 => state := s10147; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10147 => 			--6
	if (mulfprdy = '1') then state := s10148;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10147; end if;
when s10148 => state := s10149; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10149 => 			--8
	if (mulfprdy = '1') then state := s10150;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10149; end if;
when s10150 => state := s10151; 	--9
	mulfpsclr <= '0';
when s10151 => state := s10152; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10152 => 			--11
	if (mulfprdy = '1') then state := s10153;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10152; end if;
when s10153 => state := s10154; 	--12
	mulfpsclr <= '0';
when s10154 => state := s10155; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10155 => 			--14
	if (addfprdy = '1') then state := s10156;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10155; end if;
when s10156 => state := s10157; 	--15
	addfpsclr <= '0';
when s10157 => state := s10158; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10158 => 			--17
	if (addfprdy = '1') then state := s10159;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10158; end if;
when s10159 => state := s10160; 	--18
	addfpsclr <= '0';
when s10160 => state := s10161; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10161 => 			--20
	if (addfprdy = '1') then state := s10162;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10161; end if;
when s10162 => state := s10163; 	--21
	addfpsclr <= '0';
when s10163 => state := s10164; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (517, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10164 => state := s10165; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (972, 12)); -- offset LSB 924
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s10165 => state := s10166;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (973, 12)); -- offset MSB 925
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10166 => state := s10167; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10167 => 			--4
	if (fixed2floatrdy = '1') then state := s10168;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10167; end if;
when s10168 => state := s10169; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10169 => 			--6
	if (mulfprdy = '1') then state := s10170;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10169; end if;
when s10170 => state := s10171; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10171 => 			--8
	if (mulfprdy = '1') then state := s10172;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10171; end if;
when s10172 => state := s10173; 	--9
	mulfpsclr <= '0';
when s10173 => state := s10174; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10174 => 			--11
	if (mulfprdy = '1') then state := s10175;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10174; end if;
when s10175 => state := s10176; 	--12
	mulfpsclr <= '0';
when s10176 => state := s10177; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10177 => 			--14
	if (addfprdy = '1') then state := s10178;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10177; end if;
when s10178 => state := s10179; 	--15
	addfpsclr <= '0';
when s10179 => state := s10180; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10180 => 			--17
	if (addfprdy = '1') then state := s10181;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10180; end if;
when s10181 => state := s10182; 	--18
	addfpsclr <= '0';
when s10182 => state := s10183; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10183 => 			--20
	if (addfprdy = '1') then state := s10184;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10183; end if;
when s10184 => state := s10185; 	--21
	addfpsclr <= '0';
when s10185 => state := s10186; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (518, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10186 => state := s10187; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (974, 12)); -- offset LSB 926
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s10187 => state := s10188;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (975, 12)); -- offset MSB 927
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10188 => state := s10189; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10189 => 			--4
	if (fixed2floatrdy = '1') then state := s10190;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10189; end if;
when s10190 => state := s10191; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10191 => 			--6
	if (mulfprdy = '1') then state := s10192;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10191; end if;
when s10192 => state := s10193; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10193 => 			--8
	if (mulfprdy = '1') then state := s10194;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10193; end if;
when s10194 => state := s10195; 	--9
	mulfpsclr <= '0';
when s10195 => state := s10196; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10196 => 			--11
	if (mulfprdy = '1') then state := s10197;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10196; end if;
when s10197 => state := s10198; 	--12
	mulfpsclr <= '0';
when s10198 => state := s10199; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10199 => 			--14
	if (addfprdy = '1') then state := s10200;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10199; end if;
when s10200 => state := s10201; 	--15
	addfpsclr <= '0';
when s10201 => state := s10202; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10202 => 			--17
	if (addfprdy = '1') then state := s10203;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10202; end if;
when s10203 => state := s10204; 	--18
	addfpsclr <= '0';
when s10204 => state := s10205; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10205 => 			--20
	if (addfprdy = '1') then state := s10206;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10205; end if;
when s10206 => state := s10207; 	--21
	addfpsclr <= '0';
when s10207 => state := s10208; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (519, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10208 => state := s10209; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (976, 12)); -- offset LSB 928
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s10209 => state := s10210;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (977, 12)); -- offset MSB 929
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10210 => state := s10211; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10211 => 			--4
	if (fixed2floatrdy = '1') then state := s10212;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10211; end if;
when s10212 => state := s10213; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10213 => 			--6
	if (mulfprdy = '1') then state := s10214;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10213; end if;
when s10214 => state := s10215; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10215 => 			--8
	if (mulfprdy = '1') then state := s10216;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10215; end if;
when s10216 => state := s10217; 	--9
	mulfpsclr <= '0';
when s10217 => state := s10218; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10218 => 			--11
	if (mulfprdy = '1') then state := s10219;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10218; end if;
when s10219 => state := s10220; 	--12
	mulfpsclr <= '0';
when s10220 => state := s10221; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10221 => 			--14
	if (addfprdy = '1') then state := s10222;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10221; end if;
when s10222 => state := s10223; 	--15
	addfpsclr <= '0';
when s10223 => state := s10224; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10224 => 			--17
	if (addfprdy = '1') then state := s10225;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10224; end if;
when s10225 => state := s10226; 	--18
	addfpsclr <= '0';
when s10226 => state := s10227; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10227 => 			--20
	if (addfprdy = '1') then state := s10228;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10227; end if;
when s10228 => state := s10229; 	--21
	addfpsclr <= '0';
when s10229 => state := s10230; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (520, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10230 => state := s10231; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (978, 12)); -- offset LSB 930
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s10231 => state := s10232;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (979, 12)); -- offset MSB 931
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10232 => state := s10233; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10233 => 			--4
	if (fixed2floatrdy = '1') then state := s10234;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10233; end if;
when s10234 => state := s10235; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10235 => 			--6
	if (mulfprdy = '1') then state := s10236;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10235; end if;
when s10236 => state := s10237; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10237 => 			--8
	if (mulfprdy = '1') then state := s10238;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10237; end if;
when s10238 => state := s10239; 	--9
	mulfpsclr <= '0';
when s10239 => state := s10240; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10240 => 			--11
	if (mulfprdy = '1') then state := s10241;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10240; end if;
when s10241 => state := s10242; 	--12
	mulfpsclr <= '0';
when s10242 => state := s10243; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10243 => 			--14
	if (addfprdy = '1') then state := s10244;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10243; end if;
when s10244 => state := s10245; 	--15
	addfpsclr <= '0';
when s10245 => state := s10246; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10246 => 			--17
	if (addfprdy = '1') then state := s10247;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10246; end if;
when s10247 => state := s10248; 	--18
	addfpsclr <= '0';
when s10248 => state := s10249; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10249 => 			--20
	if (addfprdy = '1') then state := s10250;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10249; end if;
when s10250 => state := s10251; 	--21
	addfpsclr <= '0';
when s10251 => state := s10252; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (521, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10252 => state := s10253; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (980, 12)); -- offset LSB 932
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s10253 => state := s10254;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (981, 12)); -- offset MSB 933
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10254 => state := s10255; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10255 => 			--4
	if (fixed2floatrdy = '1') then state := s10256;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10255; end if;
when s10256 => state := s10257; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10257 => 			--6
	if (mulfprdy = '1') then state := s10258;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10257; end if;
when s10258 => state := s10259; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10259 => 			--8
	if (mulfprdy = '1') then state := s10260;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10259; end if;
when s10260 => state := s10261; 	--9
	mulfpsclr <= '0';
when s10261 => state := s10262; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10262 => 			--11
	if (mulfprdy = '1') then state := s10263;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10262; end if;
when s10263 => state := s10264; 	--12
	mulfpsclr <= '0';
when s10264 => state := s10265; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10265 => 			--14
	if (addfprdy = '1') then state := s10266;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10265; end if;
when s10266 => state := s10267; 	--15
	addfpsclr <= '0';
when s10267 => state := s10268; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10268 => 			--17
	if (addfprdy = '1') then state := s10269;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10268; end if;
when s10269 => state := s10270; 	--18
	addfpsclr <= '0';
when s10270 => state := s10271; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10271 => 			--20
	if (addfprdy = '1') then state := s10272;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10271; end if;
when s10272 => state := s10273; 	--21
	addfpsclr <= '0';
when s10273 => state := s10274; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (522, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10274 => state := s10275; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (982, 12)); -- offset LSB 934
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s10275 => state := s10276;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (983, 12)); -- offset MSB 935
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10276 => state := s10277; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10277 => 			--4
	if (fixed2floatrdy = '1') then state := s10278;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10277; end if;
when s10278 => state := s10279; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10279 => 			--6
	if (mulfprdy = '1') then state := s10280;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10279; end if;
when s10280 => state := s10281; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10281 => 			--8
	if (mulfprdy = '1') then state := s10282;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10281; end if;
when s10282 => state := s10283; 	--9
	mulfpsclr <= '0';
when s10283 => state := s10284; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10284 => 			--11
	if (mulfprdy = '1') then state := s10285;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10284; end if;
when s10285 => state := s10286; 	--12
	mulfpsclr <= '0';
when s10286 => state := s10287; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10287 => 			--14
	if (addfprdy = '1') then state := s10288;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10287; end if;
when s10288 => state := s10289; 	--15
	addfpsclr <= '0';
when s10289 => state := s10290; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10290 => 			--17
	if (addfprdy = '1') then state := s10291;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10290; end if;
when s10291 => state := s10292; 	--18
	addfpsclr <= '0';
when s10292 => state := s10293; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10293 => 			--20
	if (addfprdy = '1') then state := s10294;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10293; end if;
when s10294 => state := s10295; 	--21
	addfpsclr <= '0';
when s10295 => state := s10296; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (523, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10296 => state := s10297; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (984, 12)); -- offset LSB 936
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s10297 => state := s10298;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (985, 12)); -- offset MSB 937
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10298 => state := s10299; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10299 => 			--4
	if (fixed2floatrdy = '1') then state := s10300;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10299; end if;
when s10300 => state := s10301; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10301 => 			--6
	if (mulfprdy = '1') then state := s10302;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10301; end if;
when s10302 => state := s10303; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10303 => 			--8
	if (mulfprdy = '1') then state := s10304;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10303; end if;
when s10304 => state := s10305; 	--9
	mulfpsclr <= '0';
when s10305 => state := s10306; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10306 => 			--11
	if (mulfprdy = '1') then state := s10307;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10306; end if;
when s10307 => state := s10308; 	--12
	mulfpsclr <= '0';
when s10308 => state := s10309; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10309 => 			--14
	if (addfprdy = '1') then state := s10310;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10309; end if;
when s10310 => state := s10311; 	--15
	addfpsclr <= '0';
when s10311 => state := s10312; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10312 => 			--17
	if (addfprdy = '1') then state := s10313;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10312; end if;
when s10313 => state := s10314; 	--18
	addfpsclr <= '0';
when s10314 => state := s10315; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10315 => 			--20
	if (addfprdy = '1') then state := s10316;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10315; end if;
when s10316 => state := s10317; 	--21
	addfpsclr <= '0';
when s10317 => state := s10318; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (524, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10318 => state := s10319; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (986, 12)); -- offset LSB 938
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s10319 => state := s10320;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (987, 12)); -- offset MSB 939
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10320 => state := s10321; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10321 => 			--4
	if (fixed2floatrdy = '1') then state := s10322;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10321; end if;
when s10322 => state := s10323; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10323 => 			--6
	if (mulfprdy = '1') then state := s10324;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10323; end if;
when s10324 => state := s10325; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10325 => 			--8
	if (mulfprdy = '1') then state := s10326;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10325; end if;
when s10326 => state := s10327; 	--9
	mulfpsclr <= '0';
when s10327 => state := s10328; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10328 => 			--11
	if (mulfprdy = '1') then state := s10329;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10328; end if;
when s10329 => state := s10330; 	--12
	mulfpsclr <= '0';
when s10330 => state := s10331; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10331 => 			--14
	if (addfprdy = '1') then state := s10332;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10331; end if;
when s10332 => state := s10333; 	--15
	addfpsclr <= '0';
when s10333 => state := s10334; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10334 => 			--17
	if (addfprdy = '1') then state := s10335;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10334; end if;
when s10335 => state := s10336; 	--18
	addfpsclr <= '0';
when s10336 => state := s10337; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10337 => 			--20
	if (addfprdy = '1') then state := s10338;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10337; end if;
when s10338 => state := s10339; 	--21
	addfpsclr <= '0';
when s10339 => state := s10340; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (525, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10340 => state := s10341; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (988, 12)); -- offset LSB 940
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s10341 => state := s10342;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (989, 12)); -- offset MSB 941
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10342 => state := s10343; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10343 => 			--4
	if (fixed2floatrdy = '1') then state := s10344;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10343; end if;
when s10344 => state := s10345; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10345 => 			--6
	if (mulfprdy = '1') then state := s10346;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10345; end if;
when s10346 => state := s10347; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10347 => 			--8
	if (mulfprdy = '1') then state := s10348;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10347; end if;
when s10348 => state := s10349; 	--9
	mulfpsclr <= '0';
when s10349 => state := s10350; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10350 => 			--11
	if (mulfprdy = '1') then state := s10351;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10350; end if;
when s10351 => state := s10352; 	--12
	mulfpsclr <= '0';
when s10352 => state := s10353; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10353 => 			--14
	if (addfprdy = '1') then state := s10354;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10353; end if;
when s10354 => state := s10355; 	--15
	addfpsclr <= '0';
when s10355 => state := s10356; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10356 => 			--17
	if (addfprdy = '1') then state := s10357;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10356; end if;
when s10357 => state := s10358; 	--18
	addfpsclr <= '0';
when s10358 => state := s10359; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10359 => 			--20
	if (addfprdy = '1') then state := s10360;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10359; end if;
when s10360 => state := s10361; 	--21
	addfpsclr <= '0';
when s10361 => state := s10362; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (526, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10362 => state := s10363; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (990, 12)); -- offset LSB 942
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s10363 => state := s10364;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (991, 12)); -- offset MSB 943
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10364 => state := s10365; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10365 => 			--4
	if (fixed2floatrdy = '1') then state := s10366;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10365; end if;
when s10366 => state := s10367; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10367 => 			--6
	if (mulfprdy = '1') then state := s10368;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10367; end if;
when s10368 => state := s10369; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10369 => 			--8
	if (mulfprdy = '1') then state := s10370;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10369; end if;
when s10370 => state := s10371; 	--9
	mulfpsclr <= '0';
when s10371 => state := s10372; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10372 => 			--11
	if (mulfprdy = '1') then state := s10373;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10372; end if;
when s10373 => state := s10374; 	--12
	mulfpsclr <= '0';
when s10374 => state := s10375; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10375 => 			--14
	if (addfprdy = '1') then state := s10376;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10375; end if;
when s10376 => state := s10377; 	--15
	addfpsclr <= '0';
when s10377 => state := s10378; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10378 => 			--17
	if (addfprdy = '1') then state := s10379;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10378; end if;
when s10379 => state := s10380; 	--18
	addfpsclr <= '0';
when s10380 => state := s10381; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10381 => 			--20
	if (addfprdy = '1') then state := s10382;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10381; end if;
when s10382 => state := s10383; 	--21
	addfpsclr <= '0';
when s10383 => state := s10384; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (527, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10384 => state := s10385; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (992, 12)); -- offset LSB 944
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s10385 => state := s10386;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (993, 12)); -- offset MSB 945
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10386 => state := s10387; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10387 => 			--4
	if (fixed2floatrdy = '1') then state := s10388;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10387; end if;
when s10388 => state := s10389; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10389 => 			--6
	if (mulfprdy = '1') then state := s10390;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10389; end if;
when s10390 => state := s10391; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10391 => 			--8
	if (mulfprdy = '1') then state := s10392;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10391; end if;
when s10392 => state := s10393; 	--9
	mulfpsclr <= '0';
when s10393 => state := s10394; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10394 => 			--11
	if (mulfprdy = '1') then state := s10395;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10394; end if;
when s10395 => state := s10396; 	--12
	mulfpsclr <= '0';
when s10396 => state := s10397; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10397 => 			--14
	if (addfprdy = '1') then state := s10398;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10397; end if;
when s10398 => state := s10399; 	--15
	addfpsclr <= '0';
when s10399 => state := s10400; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10400 => 			--17
	if (addfprdy = '1') then state := s10401;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10400; end if;
when s10401 => state := s10402; 	--18
	addfpsclr <= '0';
when s10402 => state := s10403; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10403 => 			--20
	if (addfprdy = '1') then state := s10404;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10403; end if;
when s10404 => state := s10405; 	--21
	addfpsclr <= '0';
when s10405 => state := s10406; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (528, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10406 => state := s10407; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (994, 12)); -- offset LSB 946
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s10407 => state := s10408;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (995, 12)); -- offset MSB 947
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10408 => state := s10409; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10409 => 			--4
	if (fixed2floatrdy = '1') then state := s10410;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10409; end if;
when s10410 => state := s10411; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10411 => 			--6
	if (mulfprdy = '1') then state := s10412;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10411; end if;
when s10412 => state := s10413; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10413 => 			--8
	if (mulfprdy = '1') then state := s10414;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10413; end if;
when s10414 => state := s10415; 	--9
	mulfpsclr <= '0';
when s10415 => state := s10416; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10416 => 			--11
	if (mulfprdy = '1') then state := s10417;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10416; end if;
when s10417 => state := s10418; 	--12
	mulfpsclr <= '0';
when s10418 => state := s10419; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10419 => 			--14
	if (addfprdy = '1') then state := s10420;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10419; end if;
when s10420 => state := s10421; 	--15
	addfpsclr <= '0';
when s10421 => state := s10422; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10422 => 			--17
	if (addfprdy = '1') then state := s10423;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10422; end if;
when s10423 => state := s10424; 	--18
	addfpsclr <= '0';
when s10424 => state := s10425; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10425 => 			--20
	if (addfprdy = '1') then state := s10426;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10425; end if;
when s10426 => state := s10427; 	--21
	addfpsclr <= '0';
when s10427 => state := s10428; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (529, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10428 => state := s10429; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (996, 12)); -- offset LSB 948
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s10429 => state := s10430;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (997, 12)); -- offset MSB 949
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10430 => state := s10431; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10431 => 			--4
	if (fixed2floatrdy = '1') then state := s10432;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10431; end if;
when s10432 => state := s10433; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10433 => 			--6
	if (mulfprdy = '1') then state := s10434;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10433; end if;
when s10434 => state := s10435; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10435 => 			--8
	if (mulfprdy = '1') then state := s10436;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10435; end if;
when s10436 => state := s10437; 	--9
	mulfpsclr <= '0';
when s10437 => state := s10438; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10438 => 			--11
	if (mulfprdy = '1') then state := s10439;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10438; end if;
when s10439 => state := s10440; 	--12
	mulfpsclr <= '0';
when s10440 => state := s10441; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10441 => 			--14
	if (addfprdy = '1') then state := s10442;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10441; end if;
when s10442 => state := s10443; 	--15
	addfpsclr <= '0';
when s10443 => state := s10444; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10444 => 			--17
	if (addfprdy = '1') then state := s10445;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10444; end if;
when s10445 => state := s10446; 	--18
	addfpsclr <= '0';
when s10446 => state := s10447; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10447 => 			--20
	if (addfprdy = '1') then state := s10448;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10447; end if;
when s10448 => state := s10449; 	--21
	addfpsclr <= '0';
when s10449 => state := s10450; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (530, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10450 => state := s10451; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (998, 12)); -- offset LSB 950
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s10451 => state := s10452;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (999, 12)); -- offset MSB 951
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10452 => state := s10453; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10453 => 			--4
	if (fixed2floatrdy = '1') then state := s10454;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10453; end if;
when s10454 => state := s10455; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10455 => 			--6
	if (mulfprdy = '1') then state := s10456;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10455; end if;
when s10456 => state := s10457; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10457 => 			--8
	if (mulfprdy = '1') then state := s10458;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10457; end if;
when s10458 => state := s10459; 	--9
	mulfpsclr <= '0';
when s10459 => state := s10460; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10460 => 			--11
	if (mulfprdy = '1') then state := s10461;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10460; end if;
when s10461 => state := s10462; 	--12
	mulfpsclr <= '0';
when s10462 => state := s10463; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10463 => 			--14
	if (addfprdy = '1') then state := s10464;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10463; end if;
when s10464 => state := s10465; 	--15
	addfpsclr <= '0';
when s10465 => state := s10466; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10466 => 			--17
	if (addfprdy = '1') then state := s10467;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10466; end if;
when s10467 => state := s10468; 	--18
	addfpsclr <= '0';
when s10468 => state := s10469; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10469 => 			--20
	if (addfprdy = '1') then state := s10470;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10469; end if;
when s10470 => state := s10471; 	--21
	addfpsclr <= '0';
when s10471 => state := s10472; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (531, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10472 => state := s10473; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1000, 12)); -- offset LSB 952
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s10473 => state := s10474;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1001, 12)); -- offset MSB 953
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10474 => state := s10475; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10475 => 			--4
	if (fixed2floatrdy = '1') then state := s10476;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10475; end if;
when s10476 => state := s10477; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10477 => 			--6
	if (mulfprdy = '1') then state := s10478;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10477; end if;
when s10478 => state := s10479; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10479 => 			--8
	if (mulfprdy = '1') then state := s10480;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10479; end if;
when s10480 => state := s10481; 	--9
	mulfpsclr <= '0';
when s10481 => state := s10482; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10482 => 			--11
	if (mulfprdy = '1') then state := s10483;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10482; end if;
when s10483 => state := s10484; 	--12
	mulfpsclr <= '0';
when s10484 => state := s10485; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10485 => 			--14
	if (addfprdy = '1') then state := s10486;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10485; end if;
when s10486 => state := s10487; 	--15
	addfpsclr <= '0';
when s10487 => state := s10488; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10488 => 			--17
	if (addfprdy = '1') then state := s10489;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10488; end if;
when s10489 => state := s10490; 	--18
	addfpsclr <= '0';
when s10490 => state := s10491; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10491 => 			--20
	if (addfprdy = '1') then state := s10492;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10491; end if;
when s10492 => state := s10493; 	--21
	addfpsclr <= '0';
when s10493 => state := s10494; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (532, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10494 => state := s10495; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1002, 12)); -- offset LSB 954
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s10495 => state := s10496;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1003, 12)); -- offset MSB 955
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10496 => state := s10497; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10497 => 			--4
	if (fixed2floatrdy = '1') then state := s10498;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10497; end if;
when s10498 => state := s10499; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10499 => 			--6
	if (mulfprdy = '1') then state := s10500;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10499; end if;
when s10500 => state := s10501; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10501 => 			--8
	if (mulfprdy = '1') then state := s10502;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10501; end if;
when s10502 => state := s10503; 	--9
	mulfpsclr <= '0';
when s10503 => state := s10504; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10504 => 			--11
	if (mulfprdy = '1') then state := s10505;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10504; end if;
when s10505 => state := s10506; 	--12
	mulfpsclr <= '0';
when s10506 => state := s10507; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10507 => 			--14
	if (addfprdy = '1') then state := s10508;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10507; end if;
when s10508 => state := s10509; 	--15
	addfpsclr <= '0';
when s10509 => state := s10510; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10510 => 			--17
	if (addfprdy = '1') then state := s10511;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10510; end if;
when s10511 => state := s10512; 	--18
	addfpsclr <= '0';
when s10512 => state := s10513; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10513 => 			--20
	if (addfprdy = '1') then state := s10514;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10513; end if;
when s10514 => state := s10515; 	--21
	addfpsclr <= '0';
when s10515 => state := s10516; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (533, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10516 => state := s10517; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1004, 12)); -- offset LSB 956
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s10517 => state := s10518;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1005, 12)); -- offset MSB 957
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10518 => state := s10519; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10519 => 			--4
	if (fixed2floatrdy = '1') then state := s10520;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10519; end if;
when s10520 => state := s10521; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10521 => 			--6
	if (mulfprdy = '1') then state := s10522;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10521; end if;
when s10522 => state := s10523; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10523 => 			--8
	if (mulfprdy = '1') then state := s10524;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10523; end if;
when s10524 => state := s10525; 	--9
	mulfpsclr <= '0';
when s10525 => state := s10526; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10526 => 			--11
	if (mulfprdy = '1') then state := s10527;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10526; end if;
when s10527 => state := s10528; 	--12
	mulfpsclr <= '0';
when s10528 => state := s10529; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10529 => 			--14
	if (addfprdy = '1') then state := s10530;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10529; end if;
when s10530 => state := s10531; 	--15
	addfpsclr <= '0';
when s10531 => state := s10532; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10532 => 			--17
	if (addfprdy = '1') then state := s10533;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10532; end if;
when s10533 => state := s10534; 	--18
	addfpsclr <= '0';
when s10534 => state := s10535; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10535 => 			--20
	if (addfprdy = '1') then state := s10536;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10535; end if;
when s10536 => state := s10537; 	--21
	addfpsclr <= '0';
when s10537 => state := s10538; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (534, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10538 => state := s10539; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1006, 12)); -- offset LSB 958
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s10539 => state := s10540;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1007, 12)); -- offset MSB 959
	addra <= std_logic_vector (to_unsigned (14, 10)); -- OCCrowI 14
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10540 => state := s10541; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10541 => 			--4
	if (fixed2floatrdy = '1') then state := s10542;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10541; end if;
when s10542 => state := s10543; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10543 => 			--6
	if (mulfprdy = '1') then state := s10544;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10543; end if;
when s10544 => state := s10545; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10545 => 			--8
	if (mulfprdy = '1') then state := s10546;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10545; end if;
when s10546 => state := s10547; 	--9
	mulfpsclr <= '0';
when s10547 => state := s10548; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10548 => 			--11
	if (mulfprdy = '1') then state := s10549;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10548; end if;
when s10549 => state := s10550; 	--12
	mulfpsclr <= '0';
when s10550 => state := s10551; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10551 => 			--14
	if (addfprdy = '1') then state := s10552;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10551; end if;
when s10552 => state := s10553; 	--15
	addfpsclr <= '0';
when s10553 => state := s10554; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10554 => 			--17
	if (addfprdy = '1') then state := s10555;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10554; end if;
when s10555 => state := s10556; 	--18
	addfpsclr <= '0';
when s10556 => state := s10557; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10557 => 			--20
	if (addfprdy = '1') then state := s10558;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10557; end if;
when s10558 => state := s10559; 	--21
	addfpsclr <= '0';
when s10559 => state := s10560; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (535, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10560 => state := s10561; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1008, 12)); -- offset LSB 960
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s10561 => state := s10562;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1009, 12)); -- offset MSB 961
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10562 => state := s10563; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10563 => 			--4
	if (fixed2floatrdy = '1') then state := s10564;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10563; end if;
when s10564 => state := s10565; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10565 => 			--6
	if (mulfprdy = '1') then state := s10566;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10565; end if;
when s10566 => state := s10567; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10567 => 			--8
	if (mulfprdy = '1') then state := s10568;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10567; end if;
when s10568 => state := s10569; 	--9
	mulfpsclr <= '0';
when s10569 => state := s10570; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10570 => 			--11
	if (mulfprdy = '1') then state := s10571;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10570; end if;
when s10571 => state := s10572; 	--12
	mulfpsclr <= '0';
when s10572 => state := s10573; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10573 => 			--14
	if (addfprdy = '1') then state := s10574;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10573; end if;
when s10574 => state := s10575; 	--15
	addfpsclr <= '0';
when s10575 => state := s10576; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10576 => 			--17
	if (addfprdy = '1') then state := s10577;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10576; end if;
when s10577 => state := s10578; 	--18
	addfpsclr <= '0';
when s10578 => state := s10579; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10579 => 			--20
	if (addfprdy = '1') then state := s10580;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10579; end if;
when s10580 => state := s10581; 	--21
	addfpsclr <= '0';
when s10581 => state := s10582; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (536, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10582 => state := s10583; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1010, 12)); -- offset LSB 962
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s10583 => state := s10584;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1011, 12)); -- offset MSB 963
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10584 => state := s10585; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10585 => 			--4
	if (fixed2floatrdy = '1') then state := s10586;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10585; end if;
when s10586 => state := s10587; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10587 => 			--6
	if (mulfprdy = '1') then state := s10588;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10587; end if;
when s10588 => state := s10589; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10589 => 			--8
	if (mulfprdy = '1') then state := s10590;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10589; end if;
when s10590 => state := s10591; 	--9
	mulfpsclr <= '0';
when s10591 => state := s10592; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10592 => 			--11
	if (mulfprdy = '1') then state := s10593;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10592; end if;
when s10593 => state := s10594; 	--12
	mulfpsclr <= '0';
when s10594 => state := s10595; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10595 => 			--14
	if (addfprdy = '1') then state := s10596;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10595; end if;
when s10596 => state := s10597; 	--15
	addfpsclr <= '0';
when s10597 => state := s10598; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10598 => 			--17
	if (addfprdy = '1') then state := s10599;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10598; end if;
when s10599 => state := s10600; 	--18
	addfpsclr <= '0';
when s10600 => state := s10601; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10601 => 			--20
	if (addfprdy = '1') then state := s10602;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10601; end if;
when s10602 => state := s10603; 	--21
	addfpsclr <= '0';
when s10603 => state := s10604; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (537, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10604 => state := s10605; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1012, 12)); -- offset LSB 964
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s10605 => state := s10606;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1013, 12)); -- offset MSB 965
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10606 => state := s10607; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10607 => 			--4
	if (fixed2floatrdy = '1') then state := s10608;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10607; end if;
when s10608 => state := s10609; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10609 => 			--6
	if (mulfprdy = '1') then state := s10610;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10609; end if;
when s10610 => state := s10611; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10611 => 			--8
	if (mulfprdy = '1') then state := s10612;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10611; end if;
when s10612 => state := s10613; 	--9
	mulfpsclr <= '0';
when s10613 => state := s10614; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10614 => 			--11
	if (mulfprdy = '1') then state := s10615;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10614; end if;
when s10615 => state := s10616; 	--12
	mulfpsclr <= '0';
when s10616 => state := s10617; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10617 => 			--14
	if (addfprdy = '1') then state := s10618;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10617; end if;
when s10618 => state := s10619; 	--15
	addfpsclr <= '0';
when s10619 => state := s10620; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10620 => 			--17
	if (addfprdy = '1') then state := s10621;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10620; end if;
when s10621 => state := s10622; 	--18
	addfpsclr <= '0';
when s10622 => state := s10623; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10623 => 			--20
	if (addfprdy = '1') then state := s10624;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10623; end if;
when s10624 => state := s10625; 	--21
	addfpsclr <= '0';
when s10625 => state := s10626; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (538, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10626 => state := s10627; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1014, 12)); -- offset LSB 966
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s10627 => state := s10628;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1015, 12)); -- offset MSB 967
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10628 => state := s10629; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10629 => 			--4
	if (fixed2floatrdy = '1') then state := s10630;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10629; end if;
when s10630 => state := s10631; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10631 => 			--6
	if (mulfprdy = '1') then state := s10632;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10631; end if;
when s10632 => state := s10633; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10633 => 			--8
	if (mulfprdy = '1') then state := s10634;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10633; end if;
when s10634 => state := s10635; 	--9
	mulfpsclr <= '0';
when s10635 => state := s10636; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10636 => 			--11
	if (mulfprdy = '1') then state := s10637;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10636; end if;
when s10637 => state := s10638; 	--12
	mulfpsclr <= '0';
when s10638 => state := s10639; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10639 => 			--14
	if (addfprdy = '1') then state := s10640;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10639; end if;
when s10640 => state := s10641; 	--15
	addfpsclr <= '0';
when s10641 => state := s10642; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10642 => 			--17
	if (addfprdy = '1') then state := s10643;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10642; end if;
when s10643 => state := s10644; 	--18
	addfpsclr <= '0';
when s10644 => state := s10645; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10645 => 			--20
	if (addfprdy = '1') then state := s10646;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10645; end if;
when s10646 => state := s10647; 	--21
	addfpsclr <= '0';
when s10647 => state := s10648; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (539, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10648 => state := s10649; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1016, 12)); -- offset LSB 968
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s10649 => state := s10650;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1017, 12)); -- offset MSB 969
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10650 => state := s10651; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10651 => 			--4
	if (fixed2floatrdy = '1') then state := s10652;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10651; end if;
when s10652 => state := s10653; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10653 => 			--6
	if (mulfprdy = '1') then state := s10654;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10653; end if;
when s10654 => state := s10655; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10655 => 			--8
	if (mulfprdy = '1') then state := s10656;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10655; end if;
when s10656 => state := s10657; 	--9
	mulfpsclr <= '0';
when s10657 => state := s10658; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10658 => 			--11
	if (mulfprdy = '1') then state := s10659;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10658; end if;
when s10659 => state := s10660; 	--12
	mulfpsclr <= '0';
when s10660 => state := s10661; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10661 => 			--14
	if (addfprdy = '1') then state := s10662;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10661; end if;
when s10662 => state := s10663; 	--15
	addfpsclr <= '0';
when s10663 => state := s10664; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10664 => 			--17
	if (addfprdy = '1') then state := s10665;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10664; end if;
when s10665 => state := s10666; 	--18
	addfpsclr <= '0';
when s10666 => state := s10667; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10667 => 			--20
	if (addfprdy = '1') then state := s10668;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10667; end if;
when s10668 => state := s10669; 	--21
	addfpsclr <= '0';
when s10669 => state := s10670; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (540, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10670 => state := s10671; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1018, 12)); -- offset LSB 970
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s10671 => state := s10672;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1019, 12)); -- offset MSB 971
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10672 => state := s10673; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10673 => 			--4
	if (fixed2floatrdy = '1') then state := s10674;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10673; end if;
when s10674 => state := s10675; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10675 => 			--6
	if (mulfprdy = '1') then state := s10676;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10675; end if;
when s10676 => state := s10677; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10677 => 			--8
	if (mulfprdy = '1') then state := s10678;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10677; end if;
when s10678 => state := s10679; 	--9
	mulfpsclr <= '0';
when s10679 => state := s10680; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10680 => 			--11
	if (mulfprdy = '1') then state := s10681;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10680; end if;
when s10681 => state := s10682; 	--12
	mulfpsclr <= '0';
when s10682 => state := s10683; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10683 => 			--14
	if (addfprdy = '1') then state := s10684;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10683; end if;
when s10684 => state := s10685; 	--15
	addfpsclr <= '0';
when s10685 => state := s10686; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10686 => 			--17
	if (addfprdy = '1') then state := s10687;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10686; end if;
when s10687 => state := s10688; 	--18
	addfpsclr <= '0';
when s10688 => state := s10689; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10689 => 			--20
	if (addfprdy = '1') then state := s10690;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10689; end if;
when s10690 => state := s10691; 	--21
	addfpsclr <= '0';
when s10691 => state := s10692; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (541, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10692 => state := s10693; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1020, 12)); -- offset LSB 972
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s10693 => state := s10694;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1021, 12)); -- offset MSB 973
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10694 => state := s10695; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10695 => 			--4
	if (fixed2floatrdy = '1') then state := s10696;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10695; end if;
when s10696 => state := s10697; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10697 => 			--6
	if (mulfprdy = '1') then state := s10698;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10697; end if;
when s10698 => state := s10699; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10699 => 			--8
	if (mulfprdy = '1') then state := s10700;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10699; end if;
when s10700 => state := s10701; 	--9
	mulfpsclr <= '0';
when s10701 => state := s10702; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10702 => 			--11
	if (mulfprdy = '1') then state := s10703;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10702; end if;
when s10703 => state := s10704; 	--12
	mulfpsclr <= '0';
when s10704 => state := s10705; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10705 => 			--14
	if (addfprdy = '1') then state := s10706;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10705; end if;
when s10706 => state := s10707; 	--15
	addfpsclr <= '0';
when s10707 => state := s10708; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10708 => 			--17
	if (addfprdy = '1') then state := s10709;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10708; end if;
when s10709 => state := s10710; 	--18
	addfpsclr <= '0';
when s10710 => state := s10711; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10711 => 			--20
	if (addfprdy = '1') then state := s10712;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10711; end if;
when s10712 => state := s10713; 	--21
	addfpsclr <= '0';
when s10713 => state := s10714; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (542, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10714 => state := s10715; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1022, 12)); -- offset LSB 974
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s10715 => state := s10716;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1023, 12)); -- offset MSB 975
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10716 => state := s10717; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10717 => 			--4
	if (fixed2floatrdy = '1') then state := s10718;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10717; end if;
when s10718 => state := s10719; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10719 => 			--6
	if (mulfprdy = '1') then state := s10720;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10719; end if;
when s10720 => state := s10721; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10721 => 			--8
	if (mulfprdy = '1') then state := s10722;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10721; end if;
when s10722 => state := s10723; 	--9
	mulfpsclr <= '0';
when s10723 => state := s10724; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10724 => 			--11
	if (mulfprdy = '1') then state := s10725;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10724; end if;
when s10725 => state := s10726; 	--12
	mulfpsclr <= '0';
when s10726 => state := s10727; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10727 => 			--14
	if (addfprdy = '1') then state := s10728;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10727; end if;
when s10728 => state := s10729; 	--15
	addfpsclr <= '0';
when s10729 => state := s10730; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10730 => 			--17
	if (addfprdy = '1') then state := s10731;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10730; end if;
when s10731 => state := s10732; 	--18
	addfpsclr <= '0';
when s10732 => state := s10733; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10733 => 			--20
	if (addfprdy = '1') then state := s10734;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10733; end if;
when s10734 => state := s10735; 	--21
	addfpsclr <= '0';
when s10735 => state := s10736; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (543, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10736 => state := s10737; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1024, 12)); -- offset LSB 976
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s10737 => state := s10738;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1025, 12)); -- offset MSB 977
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10738 => state := s10739; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10739 => 			--4
	if (fixed2floatrdy = '1') then state := s10740;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10739; end if;
when s10740 => state := s10741; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10741 => 			--6
	if (mulfprdy = '1') then state := s10742;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10741; end if;
when s10742 => state := s10743; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10743 => 			--8
	if (mulfprdy = '1') then state := s10744;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10743; end if;
when s10744 => state := s10745; 	--9
	mulfpsclr <= '0';
when s10745 => state := s10746; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10746 => 			--11
	if (mulfprdy = '1') then state := s10747;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10746; end if;
when s10747 => state := s10748; 	--12
	mulfpsclr <= '0';
when s10748 => state := s10749; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10749 => 			--14
	if (addfprdy = '1') then state := s10750;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10749; end if;
when s10750 => state := s10751; 	--15
	addfpsclr <= '0';
when s10751 => state := s10752; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10752 => 			--17
	if (addfprdy = '1') then state := s10753;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10752; end if;
when s10753 => state := s10754; 	--18
	addfpsclr <= '0';
when s10754 => state := s10755; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10755 => 			--20
	if (addfprdy = '1') then state := s10756;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10755; end if;
when s10756 => state := s10757; 	--21
	addfpsclr <= '0';
when s10757 => state := s10758; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (544, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10758 => state := s10759; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1026, 12)); -- offset LSB 978
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s10759 => state := s10760;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1027, 12)); -- offset MSB 979
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10760 => state := s10761; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10761 => 			--4
	if (fixed2floatrdy = '1') then state := s10762;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10761; end if;
when s10762 => state := s10763; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10763 => 			--6
	if (mulfprdy = '1') then state := s10764;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10763; end if;
when s10764 => state := s10765; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10765 => 			--8
	if (mulfprdy = '1') then state := s10766;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10765; end if;
when s10766 => state := s10767; 	--9
	mulfpsclr <= '0';
when s10767 => state := s10768; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10768 => 			--11
	if (mulfprdy = '1') then state := s10769;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10768; end if;
when s10769 => state := s10770; 	--12
	mulfpsclr <= '0';
when s10770 => state := s10771; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10771 => 			--14
	if (addfprdy = '1') then state := s10772;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10771; end if;
when s10772 => state := s10773; 	--15
	addfpsclr <= '0';
when s10773 => state := s10774; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10774 => 			--17
	if (addfprdy = '1') then state := s10775;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10774; end if;
when s10775 => state := s10776; 	--18
	addfpsclr <= '0';
when s10776 => state := s10777; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10777 => 			--20
	if (addfprdy = '1') then state := s10778;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10777; end if;
when s10778 => state := s10779; 	--21
	addfpsclr <= '0';
when s10779 => state := s10780; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (545, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10780 => state := s10781; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1028, 12)); -- offset LSB 980
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s10781 => state := s10782;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1029, 12)); -- offset MSB 981
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10782 => state := s10783; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10783 => 			--4
	if (fixed2floatrdy = '1') then state := s10784;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10783; end if;
when s10784 => state := s10785; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10785 => 			--6
	if (mulfprdy = '1') then state := s10786;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10785; end if;
when s10786 => state := s10787; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10787 => 			--8
	if (mulfprdy = '1') then state := s10788;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10787; end if;
when s10788 => state := s10789; 	--9
	mulfpsclr <= '0';
when s10789 => state := s10790; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10790 => 			--11
	if (mulfprdy = '1') then state := s10791;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10790; end if;
when s10791 => state := s10792; 	--12
	mulfpsclr <= '0';
when s10792 => state := s10793; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10793 => 			--14
	if (addfprdy = '1') then state := s10794;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10793; end if;
when s10794 => state := s10795; 	--15
	addfpsclr <= '0';
when s10795 => state := s10796; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10796 => 			--17
	if (addfprdy = '1') then state := s10797;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10796; end if;
when s10797 => state := s10798; 	--18
	addfpsclr <= '0';
when s10798 => state := s10799; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10799 => 			--20
	if (addfprdy = '1') then state := s10800;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10799; end if;
when s10800 => state := s10801; 	--21
	addfpsclr <= '0';
when s10801 => state := s10802; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (546, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10802 => state := s10803; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1030, 12)); -- offset LSB 982
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s10803 => state := s10804;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1031, 12)); -- offset MSB 983
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10804 => state := s10805; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10805 => 			--4
	if (fixed2floatrdy = '1') then state := s10806;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10805; end if;
when s10806 => state := s10807; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10807 => 			--6
	if (mulfprdy = '1') then state := s10808;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10807; end if;
when s10808 => state := s10809; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10809 => 			--8
	if (mulfprdy = '1') then state := s10810;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10809; end if;
when s10810 => state := s10811; 	--9
	mulfpsclr <= '0';
when s10811 => state := s10812; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10812 => 			--11
	if (mulfprdy = '1') then state := s10813;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10812; end if;
when s10813 => state := s10814; 	--12
	mulfpsclr <= '0';
when s10814 => state := s10815; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10815 => 			--14
	if (addfprdy = '1') then state := s10816;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10815; end if;
when s10816 => state := s10817; 	--15
	addfpsclr <= '0';
when s10817 => state := s10818; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10818 => 			--17
	if (addfprdy = '1') then state := s10819;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10818; end if;
when s10819 => state := s10820; 	--18
	addfpsclr <= '0';
when s10820 => state := s10821; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10821 => 			--20
	if (addfprdy = '1') then state := s10822;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10821; end if;
when s10822 => state := s10823; 	--21
	addfpsclr <= '0';
when s10823 => state := s10824; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (547, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10824 => state := s10825; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1032, 12)); -- offset LSB 984
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s10825 => state := s10826;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1033, 12)); -- offset MSB 985
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10826 => state := s10827; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10827 => 			--4
	if (fixed2floatrdy = '1') then state := s10828;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10827; end if;
when s10828 => state := s10829; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10829 => 			--6
	if (mulfprdy = '1') then state := s10830;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10829; end if;
when s10830 => state := s10831; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10831 => 			--8
	if (mulfprdy = '1') then state := s10832;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10831; end if;
when s10832 => state := s10833; 	--9
	mulfpsclr <= '0';
when s10833 => state := s10834; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10834 => 			--11
	if (mulfprdy = '1') then state := s10835;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10834; end if;
when s10835 => state := s10836; 	--12
	mulfpsclr <= '0';
when s10836 => state := s10837; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10837 => 			--14
	if (addfprdy = '1') then state := s10838;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10837; end if;
when s10838 => state := s10839; 	--15
	addfpsclr <= '0';
when s10839 => state := s10840; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10840 => 			--17
	if (addfprdy = '1') then state := s10841;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10840; end if;
when s10841 => state := s10842; 	--18
	addfpsclr <= '0';
when s10842 => state := s10843; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10843 => 			--20
	if (addfprdy = '1') then state := s10844;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10843; end if;
when s10844 => state := s10845; 	--21
	addfpsclr <= '0';
when s10845 => state := s10846; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (548, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10846 => state := s10847; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1034, 12)); -- offset LSB 986
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s10847 => state := s10848;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1035, 12)); -- offset MSB 987
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10848 => state := s10849; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10849 => 			--4
	if (fixed2floatrdy = '1') then state := s10850;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10849; end if;
when s10850 => state := s10851; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10851 => 			--6
	if (mulfprdy = '1') then state := s10852;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10851; end if;
when s10852 => state := s10853; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10853 => 			--8
	if (mulfprdy = '1') then state := s10854;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10853; end if;
when s10854 => state := s10855; 	--9
	mulfpsclr <= '0';
when s10855 => state := s10856; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10856 => 			--11
	if (mulfprdy = '1') then state := s10857;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10856; end if;
when s10857 => state := s10858; 	--12
	mulfpsclr <= '0';
when s10858 => state := s10859; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10859 => 			--14
	if (addfprdy = '1') then state := s10860;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10859; end if;
when s10860 => state := s10861; 	--15
	addfpsclr <= '0';
when s10861 => state := s10862; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10862 => 			--17
	if (addfprdy = '1') then state := s10863;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10862; end if;
when s10863 => state := s10864; 	--18
	addfpsclr <= '0';
when s10864 => state := s10865; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10865 => 			--20
	if (addfprdy = '1') then state := s10866;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10865; end if;
when s10866 => state := s10867; 	--21
	addfpsclr <= '0';
when s10867 => state := s10868; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (549, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10868 => state := s10869; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1036, 12)); -- offset LSB 988
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s10869 => state := s10870;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1037, 12)); -- offset MSB 989
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10870 => state := s10871; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10871 => 			--4
	if (fixed2floatrdy = '1') then state := s10872;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10871; end if;
when s10872 => state := s10873; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10873 => 			--6
	if (mulfprdy = '1') then state := s10874;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10873; end if;
when s10874 => state := s10875; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10875 => 			--8
	if (mulfprdy = '1') then state := s10876;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10875; end if;
when s10876 => state := s10877; 	--9
	mulfpsclr <= '0';
when s10877 => state := s10878; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10878 => 			--11
	if (mulfprdy = '1') then state := s10879;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10878; end if;
when s10879 => state := s10880; 	--12
	mulfpsclr <= '0';
when s10880 => state := s10881; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10881 => 			--14
	if (addfprdy = '1') then state := s10882;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10881; end if;
when s10882 => state := s10883; 	--15
	addfpsclr <= '0';
when s10883 => state := s10884; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10884 => 			--17
	if (addfprdy = '1') then state := s10885;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10884; end if;
when s10885 => state := s10886; 	--18
	addfpsclr <= '0';
when s10886 => state := s10887; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10887 => 			--20
	if (addfprdy = '1') then state := s10888;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10887; end if;
when s10888 => state := s10889; 	--21
	addfpsclr <= '0';
when s10889 => state := s10890; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (550, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10890 => state := s10891; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1038, 12)); -- offset LSB 990
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s10891 => state := s10892;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1039, 12)); -- offset MSB 991
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10892 => state := s10893; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10893 => 			--4
	if (fixed2floatrdy = '1') then state := s10894;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10893; end if;
when s10894 => state := s10895; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10895 => 			--6
	if (mulfprdy = '1') then state := s10896;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10895; end if;
when s10896 => state := s10897; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10897 => 			--8
	if (mulfprdy = '1') then state := s10898;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10897; end if;
when s10898 => state := s10899; 	--9
	mulfpsclr <= '0';
when s10899 => state := s10900; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10900 => 			--11
	if (mulfprdy = '1') then state := s10901;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10900; end if;
when s10901 => state := s10902; 	--12
	mulfpsclr <= '0';
when s10902 => state := s10903; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10903 => 			--14
	if (addfprdy = '1') then state := s10904;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10903; end if;
when s10904 => state := s10905; 	--15
	addfpsclr <= '0';
when s10905 => state := s10906; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10906 => 			--17
	if (addfprdy = '1') then state := s10907;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10906; end if;
when s10907 => state := s10908; 	--18
	addfpsclr <= '0';
when s10908 => state := s10909; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10909 => 			--20
	if (addfprdy = '1') then state := s10910;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10909; end if;
when s10910 => state := s10911; 	--21
	addfpsclr <= '0';
when s10911 => state := s10912; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (551, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10912 => state := s10913; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1040, 12)); -- offset LSB 992
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s10913 => state := s10914;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1041, 12)); -- offset MSB 993
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10914 => state := s10915; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10915 => 			--4
	if (fixed2floatrdy = '1') then state := s10916;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10915; end if;
when s10916 => state := s10917; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10917 => 			--6
	if (mulfprdy = '1') then state := s10918;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10917; end if;
when s10918 => state := s10919; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10919 => 			--8
	if (mulfprdy = '1') then state := s10920;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10919; end if;
when s10920 => state := s10921; 	--9
	mulfpsclr <= '0';
when s10921 => state := s10922; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10922 => 			--11
	if (mulfprdy = '1') then state := s10923;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10922; end if;
when s10923 => state := s10924; 	--12
	mulfpsclr <= '0';
when s10924 => state := s10925; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10925 => 			--14
	if (addfprdy = '1') then state := s10926;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10925; end if;
when s10926 => state := s10927; 	--15
	addfpsclr <= '0';
when s10927 => state := s10928; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10928 => 			--17
	if (addfprdy = '1') then state := s10929;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10928; end if;
when s10929 => state := s10930; 	--18
	addfpsclr <= '0';
when s10930 => state := s10931; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10931 => 			--20
	if (addfprdy = '1') then state := s10932;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10931; end if;
when s10932 => state := s10933; 	--21
	addfpsclr <= '0';
when s10933 => state := s10934; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (552, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10934 => state := s10935; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1042, 12)); -- offset LSB 994
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s10935 => state := s10936;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1043, 12)); -- offset MSB 995
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10936 => state := s10937; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10937 => 			--4
	if (fixed2floatrdy = '1') then state := s10938;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10937; end if;
when s10938 => state := s10939; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10939 => 			--6
	if (mulfprdy = '1') then state := s10940;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10939; end if;
when s10940 => state := s10941; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10941 => 			--8
	if (mulfprdy = '1') then state := s10942;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10941; end if;
when s10942 => state := s10943; 	--9
	mulfpsclr <= '0';
when s10943 => state := s10944; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10944 => 			--11
	if (mulfprdy = '1') then state := s10945;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10944; end if;
when s10945 => state := s10946; 	--12
	mulfpsclr <= '0';
when s10946 => state := s10947; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10947 => 			--14
	if (addfprdy = '1') then state := s10948;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10947; end if;
when s10948 => state := s10949; 	--15
	addfpsclr <= '0';
when s10949 => state := s10950; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10950 => 			--17
	if (addfprdy = '1') then state := s10951;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10950; end if;
when s10951 => state := s10952; 	--18
	addfpsclr <= '0';
when s10952 => state := s10953; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10953 => 			--20
	if (addfprdy = '1') then state := s10954;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10953; end if;
when s10954 => state := s10955; 	--21
	addfpsclr <= '0';
when s10955 => state := s10956; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (553, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10956 => state := s10957; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1044, 12)); -- offset LSB 996
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s10957 => state := s10958;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1045, 12)); -- offset MSB 997
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10958 => state := s10959; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10959 => 			--4
	if (fixed2floatrdy = '1') then state := s10960;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10959; end if;
when s10960 => state := s10961; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10961 => 			--6
	if (mulfprdy = '1') then state := s10962;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10961; end if;
when s10962 => state := s10963; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10963 => 			--8
	if (mulfprdy = '1') then state := s10964;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10963; end if;
when s10964 => state := s10965; 	--9
	mulfpsclr <= '0';
when s10965 => state := s10966; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10966 => 			--11
	if (mulfprdy = '1') then state := s10967;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10966; end if;
when s10967 => state := s10968; 	--12
	mulfpsclr <= '0';
when s10968 => state := s10969; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10969 => 			--14
	if (addfprdy = '1') then state := s10970;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10969; end if;
when s10970 => state := s10971; 	--15
	addfpsclr <= '0';
when s10971 => state := s10972; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10972 => 			--17
	if (addfprdy = '1') then state := s10973;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10972; end if;
when s10973 => state := s10974; 	--18
	addfpsclr <= '0';
when s10974 => state := s10975; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10975 => 			--20
	if (addfprdy = '1') then state := s10976;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10975; end if;
when s10976 => state := s10977; 	--21
	addfpsclr <= '0';
when s10977 => state := s10978; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (554, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s10978 => state := s10979; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1046, 12)); -- offset LSB 998
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s10979 => state := s10980;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1047, 12)); -- offset MSB 999
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s10980 => state := s10981; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s10981 => 			--4
	if (fixed2floatrdy = '1') then state := s10982;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s10981; end if;
when s10982 => state := s10983; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s10983 => 			--6
	if (mulfprdy = '1') then state := s10984;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10983; end if;
when s10984 => state := s10985; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s10985 => 			--8
	if (mulfprdy = '1') then state := s10986;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10985; end if;
when s10986 => state := s10987; 	--9
	mulfpsclr <= '0';
when s10987 => state := s10988; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s10988 => 			--11
	if (mulfprdy = '1') then state := s10989;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s10988; end if;
when s10989 => state := s10990; 	--12
	mulfpsclr <= '0';
when s10990 => state := s10991; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s10991 => 			--14
	if (addfprdy = '1') then state := s10992;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10991; end if;
when s10992 => state := s10993; 	--15
	addfpsclr <= '0';
when s10993 => state := s10994; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s10994 => 			--17
	if (addfprdy = '1') then state := s10995;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10994; end if;
when s10995 => state := s10996; 	--18
	addfpsclr <= '0';
when s10996 => state := s10997; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s10997 => 			--20
	if (addfprdy = '1') then state := s10998;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s10997; end if;
when s10998 => state := s10999; 	--21
	addfpsclr <= '0';
when s10999 => state := s11000; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (555, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11000 => state := s11001; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1048, 12)); -- offset LSB 1000
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s11001 => state := s11002;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1049, 12)); -- offset MSB 1001
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11002 => state := s11003; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11003 => 			--4
	if (fixed2floatrdy = '1') then state := s11004;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11003; end if;
when s11004 => state := s11005; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11005 => 			--6
	if (mulfprdy = '1') then state := s11006;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11005; end if;
when s11006 => state := s11007; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11007 => 			--8
	if (mulfprdy = '1') then state := s11008;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11007; end if;
when s11008 => state := s11009; 	--9
	mulfpsclr <= '0';
when s11009 => state := s11010; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11010 => 			--11
	if (mulfprdy = '1') then state := s11011;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11010; end if;
when s11011 => state := s11012; 	--12
	mulfpsclr <= '0';
when s11012 => state := s11013; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11013 => 			--14
	if (addfprdy = '1') then state := s11014;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11013; end if;
when s11014 => state := s11015; 	--15
	addfpsclr <= '0';
when s11015 => state := s11016; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11016 => 			--17
	if (addfprdy = '1') then state := s11017;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11016; end if;
when s11017 => state := s11018; 	--18
	addfpsclr <= '0';
when s11018 => state := s11019; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11019 => 			--20
	if (addfprdy = '1') then state := s11020;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11019; end if;
when s11020 => state := s11021; 	--21
	addfpsclr <= '0';
when s11021 => state := s11022; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (556, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11022 => state := s11023; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1050, 12)); -- offset LSB 1002
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s11023 => state := s11024;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1051, 12)); -- offset MSB 1003
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11024 => state := s11025; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11025 => 			--4
	if (fixed2floatrdy = '1') then state := s11026;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11025; end if;
when s11026 => state := s11027; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11027 => 			--6
	if (mulfprdy = '1') then state := s11028;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11027; end if;
when s11028 => state := s11029; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11029 => 			--8
	if (mulfprdy = '1') then state := s11030;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11029; end if;
when s11030 => state := s11031; 	--9
	mulfpsclr <= '0';
when s11031 => state := s11032; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11032 => 			--11
	if (mulfprdy = '1') then state := s11033;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11032; end if;
when s11033 => state := s11034; 	--12
	mulfpsclr <= '0';
when s11034 => state := s11035; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11035 => 			--14
	if (addfprdy = '1') then state := s11036;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11035; end if;
when s11036 => state := s11037; 	--15
	addfpsclr <= '0';
when s11037 => state := s11038; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11038 => 			--17
	if (addfprdy = '1') then state := s11039;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11038; end if;
when s11039 => state := s11040; 	--18
	addfpsclr <= '0';
when s11040 => state := s11041; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11041 => 			--20
	if (addfprdy = '1') then state := s11042;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11041; end if;
when s11042 => state := s11043; 	--21
	addfpsclr <= '0';
when s11043 => state := s11044; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (557, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11044 => state := s11045; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1052, 12)); -- offset LSB 1004
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s11045 => state := s11046;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1053, 12)); -- offset MSB 1005
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11046 => state := s11047; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11047 => 			--4
	if (fixed2floatrdy = '1') then state := s11048;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11047; end if;
when s11048 => state := s11049; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11049 => 			--6
	if (mulfprdy = '1') then state := s11050;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11049; end if;
when s11050 => state := s11051; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11051 => 			--8
	if (mulfprdy = '1') then state := s11052;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11051; end if;
when s11052 => state := s11053; 	--9
	mulfpsclr <= '0';
when s11053 => state := s11054; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11054 => 			--11
	if (mulfprdy = '1') then state := s11055;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11054; end if;
when s11055 => state := s11056; 	--12
	mulfpsclr <= '0';
when s11056 => state := s11057; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11057 => 			--14
	if (addfprdy = '1') then state := s11058;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11057; end if;
when s11058 => state := s11059; 	--15
	addfpsclr <= '0';
when s11059 => state := s11060; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11060 => 			--17
	if (addfprdy = '1') then state := s11061;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11060; end if;
when s11061 => state := s11062; 	--18
	addfpsclr <= '0';
when s11062 => state := s11063; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11063 => 			--20
	if (addfprdy = '1') then state := s11064;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11063; end if;
when s11064 => state := s11065; 	--21
	addfpsclr <= '0';
when s11065 => state := s11066; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (558, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11066 => state := s11067; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1054, 12)); -- offset LSB 1006
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s11067 => state := s11068;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1055, 12)); -- offset MSB 1007
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11068 => state := s11069; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11069 => 			--4
	if (fixed2floatrdy = '1') then state := s11070;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11069; end if;
when s11070 => state := s11071; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11071 => 			--6
	if (mulfprdy = '1') then state := s11072;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11071; end if;
when s11072 => state := s11073; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11073 => 			--8
	if (mulfprdy = '1') then state := s11074;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11073; end if;
when s11074 => state := s11075; 	--9
	mulfpsclr <= '0';
when s11075 => state := s11076; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11076 => 			--11
	if (mulfprdy = '1') then state := s11077;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11076; end if;
when s11077 => state := s11078; 	--12
	mulfpsclr <= '0';
when s11078 => state := s11079; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11079 => 			--14
	if (addfprdy = '1') then state := s11080;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11079; end if;
when s11080 => state := s11081; 	--15
	addfpsclr <= '0';
when s11081 => state := s11082; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11082 => 			--17
	if (addfprdy = '1') then state := s11083;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11082; end if;
when s11083 => state := s11084; 	--18
	addfpsclr <= '0';
when s11084 => state := s11085; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11085 => 			--20
	if (addfprdy = '1') then state := s11086;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11085; end if;
when s11086 => state := s11087; 	--21
	addfpsclr <= '0';
when s11087 => state := s11088; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (559, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11088 => state := s11089; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1056, 12)); -- offset LSB 1008
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s11089 => state := s11090;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1057, 12)); -- offset MSB 1009
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11090 => state := s11091; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11091 => 			--4
	if (fixed2floatrdy = '1') then state := s11092;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11091; end if;
when s11092 => state := s11093; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11093 => 			--6
	if (mulfprdy = '1') then state := s11094;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11093; end if;
when s11094 => state := s11095; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11095 => 			--8
	if (mulfprdy = '1') then state := s11096;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11095; end if;
when s11096 => state := s11097; 	--9
	mulfpsclr <= '0';
when s11097 => state := s11098; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11098 => 			--11
	if (mulfprdy = '1') then state := s11099;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11098; end if;
when s11099 => state := s11100; 	--12
	mulfpsclr <= '0';
when s11100 => state := s11101; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11101 => 			--14
	if (addfprdy = '1') then state := s11102;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11101; end if;
when s11102 => state := s11103; 	--15
	addfpsclr <= '0';
when s11103 => state := s11104; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11104 => 			--17
	if (addfprdy = '1') then state := s11105;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11104; end if;
when s11105 => state := s11106; 	--18
	addfpsclr <= '0';
when s11106 => state := s11107; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11107 => 			--20
	if (addfprdy = '1') then state := s11108;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11107; end if;
when s11108 => state := s11109; 	--21
	addfpsclr <= '0';
when s11109 => state := s11110; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (560, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11110 => state := s11111; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1058, 12)); -- offset LSB 1010
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s11111 => state := s11112;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1059, 12)); -- offset MSB 1011
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11112 => state := s11113; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11113 => 			--4
	if (fixed2floatrdy = '1') then state := s11114;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11113; end if;
when s11114 => state := s11115; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11115 => 			--6
	if (mulfprdy = '1') then state := s11116;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11115; end if;
when s11116 => state := s11117; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11117 => 			--8
	if (mulfprdy = '1') then state := s11118;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11117; end if;
when s11118 => state := s11119; 	--9
	mulfpsclr <= '0';
when s11119 => state := s11120; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11120 => 			--11
	if (mulfprdy = '1') then state := s11121;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11120; end if;
when s11121 => state := s11122; 	--12
	mulfpsclr <= '0';
when s11122 => state := s11123; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11123 => 			--14
	if (addfprdy = '1') then state := s11124;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11123; end if;
when s11124 => state := s11125; 	--15
	addfpsclr <= '0';
when s11125 => state := s11126; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11126 => 			--17
	if (addfprdy = '1') then state := s11127;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11126; end if;
when s11127 => state := s11128; 	--18
	addfpsclr <= '0';
when s11128 => state := s11129; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11129 => 			--20
	if (addfprdy = '1') then state := s11130;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11129; end if;
when s11130 => state := s11131; 	--21
	addfpsclr <= '0';
when s11131 => state := s11132; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (561, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11132 => state := s11133; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1060, 12)); -- offset LSB 1012
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s11133 => state := s11134;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1061, 12)); -- offset MSB 1013
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11134 => state := s11135; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11135 => 			--4
	if (fixed2floatrdy = '1') then state := s11136;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11135; end if;
when s11136 => state := s11137; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11137 => 			--6
	if (mulfprdy = '1') then state := s11138;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11137; end if;
when s11138 => state := s11139; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11139 => 			--8
	if (mulfprdy = '1') then state := s11140;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11139; end if;
when s11140 => state := s11141; 	--9
	mulfpsclr <= '0';
when s11141 => state := s11142; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11142 => 			--11
	if (mulfprdy = '1') then state := s11143;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11142; end if;
when s11143 => state := s11144; 	--12
	mulfpsclr <= '0';
when s11144 => state := s11145; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11145 => 			--14
	if (addfprdy = '1') then state := s11146;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11145; end if;
when s11146 => state := s11147; 	--15
	addfpsclr <= '0';
when s11147 => state := s11148; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11148 => 			--17
	if (addfprdy = '1') then state := s11149;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11148; end if;
when s11149 => state := s11150; 	--18
	addfpsclr <= '0';
when s11150 => state := s11151; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11151 => 			--20
	if (addfprdy = '1') then state := s11152;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11151; end if;
when s11152 => state := s11153; 	--21
	addfpsclr <= '0';
when s11153 => state := s11154; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (562, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11154 => state := s11155; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1062, 12)); -- offset LSB 1014
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s11155 => state := s11156;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1063, 12)); -- offset MSB 1015
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11156 => state := s11157; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11157 => 			--4
	if (fixed2floatrdy = '1') then state := s11158;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11157; end if;
when s11158 => state := s11159; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11159 => 			--6
	if (mulfprdy = '1') then state := s11160;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11159; end if;
when s11160 => state := s11161; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11161 => 			--8
	if (mulfprdy = '1') then state := s11162;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11161; end if;
when s11162 => state := s11163; 	--9
	mulfpsclr <= '0';
when s11163 => state := s11164; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11164 => 			--11
	if (mulfprdy = '1') then state := s11165;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11164; end if;
when s11165 => state := s11166; 	--12
	mulfpsclr <= '0';
when s11166 => state := s11167; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11167 => 			--14
	if (addfprdy = '1') then state := s11168;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11167; end if;
when s11168 => state := s11169; 	--15
	addfpsclr <= '0';
when s11169 => state := s11170; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11170 => 			--17
	if (addfprdy = '1') then state := s11171;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11170; end if;
when s11171 => state := s11172; 	--18
	addfpsclr <= '0';
when s11172 => state := s11173; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11173 => 			--20
	if (addfprdy = '1') then state := s11174;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11173; end if;
when s11174 => state := s11175; 	--21
	addfpsclr <= '0';
when s11175 => state := s11176; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (563, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11176 => state := s11177; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1064, 12)); -- offset LSB 1016
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s11177 => state := s11178;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1065, 12)); -- offset MSB 1017
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11178 => state := s11179; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11179 => 			--4
	if (fixed2floatrdy = '1') then state := s11180;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11179; end if;
when s11180 => state := s11181; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11181 => 			--6
	if (mulfprdy = '1') then state := s11182;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11181; end if;
when s11182 => state := s11183; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11183 => 			--8
	if (mulfprdy = '1') then state := s11184;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11183; end if;
when s11184 => state := s11185; 	--9
	mulfpsclr <= '0';
when s11185 => state := s11186; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11186 => 			--11
	if (mulfprdy = '1') then state := s11187;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11186; end if;
when s11187 => state := s11188; 	--12
	mulfpsclr <= '0';
when s11188 => state := s11189; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11189 => 			--14
	if (addfprdy = '1') then state := s11190;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11189; end if;
when s11190 => state := s11191; 	--15
	addfpsclr <= '0';
when s11191 => state := s11192; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11192 => 			--17
	if (addfprdy = '1') then state := s11193;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11192; end if;
when s11193 => state := s11194; 	--18
	addfpsclr <= '0';
when s11194 => state := s11195; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11195 => 			--20
	if (addfprdy = '1') then state := s11196;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11195; end if;
when s11196 => state := s11197; 	--21
	addfpsclr <= '0';
when s11197 => state := s11198; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (564, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11198 => state := s11199; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1066, 12)); -- offset LSB 1018
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s11199 => state := s11200;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1067, 12)); -- offset MSB 1019
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11200 => state := s11201; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11201 => 			--4
	if (fixed2floatrdy = '1') then state := s11202;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11201; end if;
when s11202 => state := s11203; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11203 => 			--6
	if (mulfprdy = '1') then state := s11204;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11203; end if;
when s11204 => state := s11205; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11205 => 			--8
	if (mulfprdy = '1') then state := s11206;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11205; end if;
when s11206 => state := s11207; 	--9
	mulfpsclr <= '0';
when s11207 => state := s11208; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11208 => 			--11
	if (mulfprdy = '1') then state := s11209;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11208; end if;
when s11209 => state := s11210; 	--12
	mulfpsclr <= '0';
when s11210 => state := s11211; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11211 => 			--14
	if (addfprdy = '1') then state := s11212;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11211; end if;
when s11212 => state := s11213; 	--15
	addfpsclr <= '0';
when s11213 => state := s11214; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11214 => 			--17
	if (addfprdy = '1') then state := s11215;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11214; end if;
when s11215 => state := s11216; 	--18
	addfpsclr <= '0';
when s11216 => state := s11217; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11217 => 			--20
	if (addfprdy = '1') then state := s11218;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11217; end if;
when s11218 => state := s11219; 	--21
	addfpsclr <= '0';
when s11219 => state := s11220; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (565, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11220 => state := s11221; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1068, 12)); -- offset LSB 1020
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s11221 => state := s11222;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1069, 12)); -- offset MSB 1021
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11222 => state := s11223; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11223 => 			--4
	if (fixed2floatrdy = '1') then state := s11224;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11223; end if;
when s11224 => state := s11225; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11225 => 			--6
	if (mulfprdy = '1') then state := s11226;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11225; end if;
when s11226 => state := s11227; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11227 => 			--8
	if (mulfprdy = '1') then state := s11228;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11227; end if;
when s11228 => state := s11229; 	--9
	mulfpsclr <= '0';
when s11229 => state := s11230; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11230 => 			--11
	if (mulfprdy = '1') then state := s11231;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11230; end if;
when s11231 => state := s11232; 	--12
	mulfpsclr <= '0';
when s11232 => state := s11233; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11233 => 			--14
	if (addfprdy = '1') then state := s11234;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11233; end if;
when s11234 => state := s11235; 	--15
	addfpsclr <= '0';
when s11235 => state := s11236; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11236 => 			--17
	if (addfprdy = '1') then state := s11237;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11236; end if;
when s11237 => state := s11238; 	--18
	addfpsclr <= '0';
when s11238 => state := s11239; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11239 => 			--20
	if (addfprdy = '1') then state := s11240;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11239; end if;
when s11240 => state := s11241; 	--21
	addfpsclr <= '0';
when s11241 => state := s11242; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (566, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11242 => state := s11243; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1070, 12)); -- offset LSB 1022
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s11243 => state := s11244;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1071, 12)); -- offset MSB 1023
	addra <= std_logic_vector (to_unsigned (15, 10)); -- OCCrowI 15
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11244 => state := s11245; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11245 => 			--4
	if (fixed2floatrdy = '1') then state := s11246;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11245; end if;
when s11246 => state := s11247; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11247 => 			--6
	if (mulfprdy = '1') then state := s11248;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11247; end if;
when s11248 => state := s11249; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11249 => 			--8
	if (mulfprdy = '1') then state := s11250;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11249; end if;
when s11250 => state := s11251; 	--9
	mulfpsclr <= '0';
when s11251 => state := s11252; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11252 => 			--11
	if (mulfprdy = '1') then state := s11253;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11252; end if;
when s11253 => state := s11254; 	--12
	mulfpsclr <= '0';
when s11254 => state := s11255; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11255 => 			--14
	if (addfprdy = '1') then state := s11256;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11255; end if;
when s11256 => state := s11257; 	--15
	addfpsclr <= '0';
when s11257 => state := s11258; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11258 => 			--17
	if (addfprdy = '1') then state := s11259;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11258; end if;
when s11259 => state := s11260; 	--18
	addfpsclr <= '0';
when s11260 => state := s11261; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11261 => 			--20
	if (addfprdy = '1') then state := s11262;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11261; end if;
when s11262 => state := s11263; 	--21
	addfpsclr <= '0';
when s11263 => state := s11264; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (567, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11264 => state := s11265; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1072, 12)); -- offset LSB 1024
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s11265 => state := s11266;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1073, 12)); -- offset MSB 1025
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11266 => state := s11267; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11267 => 			--4
	if (fixed2floatrdy = '1') then state := s11268;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11267; end if;
when s11268 => state := s11269; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11269 => 			--6
	if (mulfprdy = '1') then state := s11270;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11269; end if;
when s11270 => state := s11271; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11271 => 			--8
	if (mulfprdy = '1') then state := s11272;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11271; end if;
when s11272 => state := s11273; 	--9
	mulfpsclr <= '0';
when s11273 => state := s11274; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11274 => 			--11
	if (mulfprdy = '1') then state := s11275;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11274; end if;
when s11275 => state := s11276; 	--12
	mulfpsclr <= '0';
when s11276 => state := s11277; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11277 => 			--14
	if (addfprdy = '1') then state := s11278;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11277; end if;
when s11278 => state := s11279; 	--15
	addfpsclr <= '0';
when s11279 => state := s11280; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11280 => 			--17
	if (addfprdy = '1') then state := s11281;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11280; end if;
when s11281 => state := s11282; 	--18
	addfpsclr <= '0';
when s11282 => state := s11283; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11283 => 			--20
	if (addfprdy = '1') then state := s11284;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11283; end if;
when s11284 => state := s11285; 	--21
	addfpsclr <= '0';
when s11285 => state := s11286; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (568, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11286 => state := s11287; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1074, 12)); -- offset LSB 1026
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s11287 => state := s11288;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1075, 12)); -- offset MSB 1027
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11288 => state := s11289; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11289 => 			--4
	if (fixed2floatrdy = '1') then state := s11290;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11289; end if;
when s11290 => state := s11291; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11291 => 			--6
	if (mulfprdy = '1') then state := s11292;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11291; end if;
when s11292 => state := s11293; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11293 => 			--8
	if (mulfprdy = '1') then state := s11294;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11293; end if;
when s11294 => state := s11295; 	--9
	mulfpsclr <= '0';
when s11295 => state := s11296; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11296 => 			--11
	if (mulfprdy = '1') then state := s11297;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11296; end if;
when s11297 => state := s11298; 	--12
	mulfpsclr <= '0';
when s11298 => state := s11299; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11299 => 			--14
	if (addfprdy = '1') then state := s11300;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11299; end if;
when s11300 => state := s11301; 	--15
	addfpsclr <= '0';
when s11301 => state := s11302; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11302 => 			--17
	if (addfprdy = '1') then state := s11303;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11302; end if;
when s11303 => state := s11304; 	--18
	addfpsclr <= '0';
when s11304 => state := s11305; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11305 => 			--20
	if (addfprdy = '1') then state := s11306;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11305; end if;
when s11306 => state := s11307; 	--21
	addfpsclr <= '0';
when s11307 => state := s11308; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (569, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11308 => state := s11309; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1076, 12)); -- offset LSB 1028
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s11309 => state := s11310;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1077, 12)); -- offset MSB 1029
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11310 => state := s11311; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11311 => 			--4
	if (fixed2floatrdy = '1') then state := s11312;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11311; end if;
when s11312 => state := s11313; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11313 => 			--6
	if (mulfprdy = '1') then state := s11314;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11313; end if;
when s11314 => state := s11315; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11315 => 			--8
	if (mulfprdy = '1') then state := s11316;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11315; end if;
when s11316 => state := s11317; 	--9
	mulfpsclr <= '0';
when s11317 => state := s11318; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11318 => 			--11
	if (mulfprdy = '1') then state := s11319;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11318; end if;
when s11319 => state := s11320; 	--12
	mulfpsclr <= '0';
when s11320 => state := s11321; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11321 => 			--14
	if (addfprdy = '1') then state := s11322;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11321; end if;
when s11322 => state := s11323; 	--15
	addfpsclr <= '0';
when s11323 => state := s11324; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11324 => 			--17
	if (addfprdy = '1') then state := s11325;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11324; end if;
when s11325 => state := s11326; 	--18
	addfpsclr <= '0';
when s11326 => state := s11327; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11327 => 			--20
	if (addfprdy = '1') then state := s11328;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11327; end if;
when s11328 => state := s11329; 	--21
	addfpsclr <= '0';
when s11329 => state := s11330; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (570, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11330 => state := s11331; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1078, 12)); -- offset LSB 1030
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s11331 => state := s11332;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1079, 12)); -- offset MSB 1031
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11332 => state := s11333; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11333 => 			--4
	if (fixed2floatrdy = '1') then state := s11334;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11333; end if;
when s11334 => state := s11335; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11335 => 			--6
	if (mulfprdy = '1') then state := s11336;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11335; end if;
when s11336 => state := s11337; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11337 => 			--8
	if (mulfprdy = '1') then state := s11338;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11337; end if;
when s11338 => state := s11339; 	--9
	mulfpsclr <= '0';
when s11339 => state := s11340; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11340 => 			--11
	if (mulfprdy = '1') then state := s11341;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11340; end if;
when s11341 => state := s11342; 	--12
	mulfpsclr <= '0';
when s11342 => state := s11343; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11343 => 			--14
	if (addfprdy = '1') then state := s11344;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11343; end if;
when s11344 => state := s11345; 	--15
	addfpsclr <= '0';
when s11345 => state := s11346; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11346 => 			--17
	if (addfprdy = '1') then state := s11347;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11346; end if;
when s11347 => state := s11348; 	--18
	addfpsclr <= '0';
when s11348 => state := s11349; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11349 => 			--20
	if (addfprdy = '1') then state := s11350;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11349; end if;
when s11350 => state := s11351; 	--21
	addfpsclr <= '0';
when s11351 => state := s11352; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (571, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11352 => state := s11353; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1080, 12)); -- offset LSB 1032
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s11353 => state := s11354;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1081, 12)); -- offset MSB 1033
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11354 => state := s11355; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11355 => 			--4
	if (fixed2floatrdy = '1') then state := s11356;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11355; end if;
when s11356 => state := s11357; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11357 => 			--6
	if (mulfprdy = '1') then state := s11358;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11357; end if;
when s11358 => state := s11359; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11359 => 			--8
	if (mulfprdy = '1') then state := s11360;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11359; end if;
when s11360 => state := s11361; 	--9
	mulfpsclr <= '0';
when s11361 => state := s11362; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11362 => 			--11
	if (mulfprdy = '1') then state := s11363;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11362; end if;
when s11363 => state := s11364; 	--12
	mulfpsclr <= '0';
when s11364 => state := s11365; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11365 => 			--14
	if (addfprdy = '1') then state := s11366;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11365; end if;
when s11366 => state := s11367; 	--15
	addfpsclr <= '0';
when s11367 => state := s11368; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11368 => 			--17
	if (addfprdy = '1') then state := s11369;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11368; end if;
when s11369 => state := s11370; 	--18
	addfpsclr <= '0';
when s11370 => state := s11371; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11371 => 			--20
	if (addfprdy = '1') then state := s11372;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11371; end if;
when s11372 => state := s11373; 	--21
	addfpsclr <= '0';
when s11373 => state := s11374; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (572, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11374 => state := s11375; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1082, 12)); -- offset LSB 1034
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s11375 => state := s11376;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1083, 12)); -- offset MSB 1035
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11376 => state := s11377; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11377 => 			--4
	if (fixed2floatrdy = '1') then state := s11378;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11377; end if;
when s11378 => state := s11379; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11379 => 			--6
	if (mulfprdy = '1') then state := s11380;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11379; end if;
when s11380 => state := s11381; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11381 => 			--8
	if (mulfprdy = '1') then state := s11382;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11381; end if;
when s11382 => state := s11383; 	--9
	mulfpsclr <= '0';
when s11383 => state := s11384; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11384 => 			--11
	if (mulfprdy = '1') then state := s11385;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11384; end if;
when s11385 => state := s11386; 	--12
	mulfpsclr <= '0';
when s11386 => state := s11387; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11387 => 			--14
	if (addfprdy = '1') then state := s11388;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11387; end if;
when s11388 => state := s11389; 	--15
	addfpsclr <= '0';
when s11389 => state := s11390; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11390 => 			--17
	if (addfprdy = '1') then state := s11391;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11390; end if;
when s11391 => state := s11392; 	--18
	addfpsclr <= '0';
when s11392 => state := s11393; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11393 => 			--20
	if (addfprdy = '1') then state := s11394;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11393; end if;
when s11394 => state := s11395; 	--21
	addfpsclr <= '0';
when s11395 => state := s11396; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (573, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11396 => state := s11397; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1084, 12)); -- offset LSB 1036
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s11397 => state := s11398;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1085, 12)); -- offset MSB 1037
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11398 => state := s11399; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11399 => 			--4
	if (fixed2floatrdy = '1') then state := s11400;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11399; end if;
when s11400 => state := s11401; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11401 => 			--6
	if (mulfprdy = '1') then state := s11402;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11401; end if;
when s11402 => state := s11403; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11403 => 			--8
	if (mulfprdy = '1') then state := s11404;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11403; end if;
when s11404 => state := s11405; 	--9
	mulfpsclr <= '0';
when s11405 => state := s11406; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11406 => 			--11
	if (mulfprdy = '1') then state := s11407;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11406; end if;
when s11407 => state := s11408; 	--12
	mulfpsclr <= '0';
when s11408 => state := s11409; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11409 => 			--14
	if (addfprdy = '1') then state := s11410;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11409; end if;
when s11410 => state := s11411; 	--15
	addfpsclr <= '0';
when s11411 => state := s11412; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11412 => 			--17
	if (addfprdy = '1') then state := s11413;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11412; end if;
when s11413 => state := s11414; 	--18
	addfpsclr <= '0';
when s11414 => state := s11415; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11415 => 			--20
	if (addfprdy = '1') then state := s11416;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11415; end if;
when s11416 => state := s11417; 	--21
	addfpsclr <= '0';
when s11417 => state := s11418; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (574, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11418 => state := s11419; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1086, 12)); -- offset LSB 1038
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s11419 => state := s11420;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1087, 12)); -- offset MSB 1039
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11420 => state := s11421; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11421 => 			--4
	if (fixed2floatrdy = '1') then state := s11422;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11421; end if;
when s11422 => state := s11423; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11423 => 			--6
	if (mulfprdy = '1') then state := s11424;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11423; end if;
when s11424 => state := s11425; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11425 => 			--8
	if (mulfprdy = '1') then state := s11426;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11425; end if;
when s11426 => state := s11427; 	--9
	mulfpsclr <= '0';
when s11427 => state := s11428; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11428 => 			--11
	if (mulfprdy = '1') then state := s11429;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11428; end if;
when s11429 => state := s11430; 	--12
	mulfpsclr <= '0';
when s11430 => state := s11431; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11431 => 			--14
	if (addfprdy = '1') then state := s11432;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11431; end if;
when s11432 => state := s11433; 	--15
	addfpsclr <= '0';
when s11433 => state := s11434; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11434 => 			--17
	if (addfprdy = '1') then state := s11435;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11434; end if;
when s11435 => state := s11436; 	--18
	addfpsclr <= '0';
when s11436 => state := s11437; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11437 => 			--20
	if (addfprdy = '1') then state := s11438;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11437; end if;
when s11438 => state := s11439; 	--21
	addfpsclr <= '0';
when s11439 => state := s11440; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (575, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11440 => state := s11441; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1088, 12)); -- offset LSB 1040
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s11441 => state := s11442;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1089, 12)); -- offset MSB 1041
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11442 => state := s11443; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11443 => 			--4
	if (fixed2floatrdy = '1') then state := s11444;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11443; end if;
when s11444 => state := s11445; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11445 => 			--6
	if (mulfprdy = '1') then state := s11446;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11445; end if;
when s11446 => state := s11447; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11447 => 			--8
	if (mulfprdy = '1') then state := s11448;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11447; end if;
when s11448 => state := s11449; 	--9
	mulfpsclr <= '0';
when s11449 => state := s11450; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11450 => 			--11
	if (mulfprdy = '1') then state := s11451;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11450; end if;
when s11451 => state := s11452; 	--12
	mulfpsclr <= '0';
when s11452 => state := s11453; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11453 => 			--14
	if (addfprdy = '1') then state := s11454;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11453; end if;
when s11454 => state := s11455; 	--15
	addfpsclr <= '0';
when s11455 => state := s11456; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11456 => 			--17
	if (addfprdy = '1') then state := s11457;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11456; end if;
when s11457 => state := s11458; 	--18
	addfpsclr <= '0';
when s11458 => state := s11459; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11459 => 			--20
	if (addfprdy = '1') then state := s11460;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11459; end if;
when s11460 => state := s11461; 	--21
	addfpsclr <= '0';
when s11461 => state := s11462; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (576, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11462 => state := s11463; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1090, 12)); -- offset LSB 1042
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s11463 => state := s11464;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1091, 12)); -- offset MSB 1043
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11464 => state := s11465; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11465 => 			--4
	if (fixed2floatrdy = '1') then state := s11466;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11465; end if;
when s11466 => state := s11467; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11467 => 			--6
	if (mulfprdy = '1') then state := s11468;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11467; end if;
when s11468 => state := s11469; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11469 => 			--8
	if (mulfprdy = '1') then state := s11470;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11469; end if;
when s11470 => state := s11471; 	--9
	mulfpsclr <= '0';
when s11471 => state := s11472; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11472 => 			--11
	if (mulfprdy = '1') then state := s11473;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11472; end if;
when s11473 => state := s11474; 	--12
	mulfpsclr <= '0';
when s11474 => state := s11475; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11475 => 			--14
	if (addfprdy = '1') then state := s11476;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11475; end if;
when s11476 => state := s11477; 	--15
	addfpsclr <= '0';
when s11477 => state := s11478; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11478 => 			--17
	if (addfprdy = '1') then state := s11479;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11478; end if;
when s11479 => state := s11480; 	--18
	addfpsclr <= '0';
when s11480 => state := s11481; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11481 => 			--20
	if (addfprdy = '1') then state := s11482;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11481; end if;
when s11482 => state := s11483; 	--21
	addfpsclr <= '0';
when s11483 => state := s11484; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (577, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11484 => state := s11485; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1092, 12)); -- offset LSB 1044
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s11485 => state := s11486;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1093, 12)); -- offset MSB 1045
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11486 => state := s11487; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11487 => 			--4
	if (fixed2floatrdy = '1') then state := s11488;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11487; end if;
when s11488 => state := s11489; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11489 => 			--6
	if (mulfprdy = '1') then state := s11490;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11489; end if;
when s11490 => state := s11491; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11491 => 			--8
	if (mulfprdy = '1') then state := s11492;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11491; end if;
when s11492 => state := s11493; 	--9
	mulfpsclr <= '0';
when s11493 => state := s11494; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11494 => 			--11
	if (mulfprdy = '1') then state := s11495;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11494; end if;
when s11495 => state := s11496; 	--12
	mulfpsclr <= '0';
when s11496 => state := s11497; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11497 => 			--14
	if (addfprdy = '1') then state := s11498;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11497; end if;
when s11498 => state := s11499; 	--15
	addfpsclr <= '0';
when s11499 => state := s11500; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11500 => 			--17
	if (addfprdy = '1') then state := s11501;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11500; end if;
when s11501 => state := s11502; 	--18
	addfpsclr <= '0';
when s11502 => state := s11503; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11503 => 			--20
	if (addfprdy = '1') then state := s11504;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11503; end if;
when s11504 => state := s11505; 	--21
	addfpsclr <= '0';
when s11505 => state := s11506; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (578, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11506 => state := s11507; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1094, 12)); -- offset LSB 1046
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s11507 => state := s11508;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1095, 12)); -- offset MSB 1047
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11508 => state := s11509; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11509 => 			--4
	if (fixed2floatrdy = '1') then state := s11510;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11509; end if;
when s11510 => state := s11511; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11511 => 			--6
	if (mulfprdy = '1') then state := s11512;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11511; end if;
when s11512 => state := s11513; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11513 => 			--8
	if (mulfprdy = '1') then state := s11514;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11513; end if;
when s11514 => state := s11515; 	--9
	mulfpsclr <= '0';
when s11515 => state := s11516; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11516 => 			--11
	if (mulfprdy = '1') then state := s11517;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11516; end if;
when s11517 => state := s11518; 	--12
	mulfpsclr <= '0';
when s11518 => state := s11519; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11519 => 			--14
	if (addfprdy = '1') then state := s11520;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11519; end if;
when s11520 => state := s11521; 	--15
	addfpsclr <= '0';
when s11521 => state := s11522; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11522 => 			--17
	if (addfprdy = '1') then state := s11523;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11522; end if;
when s11523 => state := s11524; 	--18
	addfpsclr <= '0';
when s11524 => state := s11525; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11525 => 			--20
	if (addfprdy = '1') then state := s11526;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11525; end if;
when s11526 => state := s11527; 	--21
	addfpsclr <= '0';
when s11527 => state := s11528; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (579, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11528 => state := s11529; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1096, 12)); -- offset LSB 1048
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s11529 => state := s11530;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1097, 12)); -- offset MSB 1049
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11530 => state := s11531; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11531 => 			--4
	if (fixed2floatrdy = '1') then state := s11532;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11531; end if;
when s11532 => state := s11533; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11533 => 			--6
	if (mulfprdy = '1') then state := s11534;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11533; end if;
when s11534 => state := s11535; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11535 => 			--8
	if (mulfprdy = '1') then state := s11536;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11535; end if;
when s11536 => state := s11537; 	--9
	mulfpsclr <= '0';
when s11537 => state := s11538; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11538 => 			--11
	if (mulfprdy = '1') then state := s11539;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11538; end if;
when s11539 => state := s11540; 	--12
	mulfpsclr <= '0';
when s11540 => state := s11541; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11541 => 			--14
	if (addfprdy = '1') then state := s11542;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11541; end if;
when s11542 => state := s11543; 	--15
	addfpsclr <= '0';
when s11543 => state := s11544; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11544 => 			--17
	if (addfprdy = '1') then state := s11545;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11544; end if;
when s11545 => state := s11546; 	--18
	addfpsclr <= '0';
when s11546 => state := s11547; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11547 => 			--20
	if (addfprdy = '1') then state := s11548;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11547; end if;
when s11548 => state := s11549; 	--21
	addfpsclr <= '0';
when s11549 => state := s11550; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (580, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11550 => state := s11551; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1098, 12)); -- offset LSB 1050
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s11551 => state := s11552;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1099, 12)); -- offset MSB 1051
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11552 => state := s11553; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11553 => 			--4
	if (fixed2floatrdy = '1') then state := s11554;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11553; end if;
when s11554 => state := s11555; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11555 => 			--6
	if (mulfprdy = '1') then state := s11556;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11555; end if;
when s11556 => state := s11557; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11557 => 			--8
	if (mulfprdy = '1') then state := s11558;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11557; end if;
when s11558 => state := s11559; 	--9
	mulfpsclr <= '0';
when s11559 => state := s11560; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11560 => 			--11
	if (mulfprdy = '1') then state := s11561;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11560; end if;
when s11561 => state := s11562; 	--12
	mulfpsclr <= '0';
when s11562 => state := s11563; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11563 => 			--14
	if (addfprdy = '1') then state := s11564;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11563; end if;
when s11564 => state := s11565; 	--15
	addfpsclr <= '0';
when s11565 => state := s11566; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11566 => 			--17
	if (addfprdy = '1') then state := s11567;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11566; end if;
when s11567 => state := s11568; 	--18
	addfpsclr <= '0';
when s11568 => state := s11569; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11569 => 			--20
	if (addfprdy = '1') then state := s11570;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11569; end if;
when s11570 => state := s11571; 	--21
	addfpsclr <= '0';
when s11571 => state := s11572; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (581, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11572 => state := s11573; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1100, 12)); -- offset LSB 1052
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s11573 => state := s11574;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1101, 12)); -- offset MSB 1053
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11574 => state := s11575; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11575 => 			--4
	if (fixed2floatrdy = '1') then state := s11576;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11575; end if;
when s11576 => state := s11577; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11577 => 			--6
	if (mulfprdy = '1') then state := s11578;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11577; end if;
when s11578 => state := s11579; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11579 => 			--8
	if (mulfprdy = '1') then state := s11580;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11579; end if;
when s11580 => state := s11581; 	--9
	mulfpsclr <= '0';
when s11581 => state := s11582; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11582 => 			--11
	if (mulfprdy = '1') then state := s11583;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11582; end if;
when s11583 => state := s11584; 	--12
	mulfpsclr <= '0';
when s11584 => state := s11585; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11585 => 			--14
	if (addfprdy = '1') then state := s11586;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11585; end if;
when s11586 => state := s11587; 	--15
	addfpsclr <= '0';
when s11587 => state := s11588; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11588 => 			--17
	if (addfprdy = '1') then state := s11589;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11588; end if;
when s11589 => state := s11590; 	--18
	addfpsclr <= '0';
when s11590 => state := s11591; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11591 => 			--20
	if (addfprdy = '1') then state := s11592;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11591; end if;
when s11592 => state := s11593; 	--21
	addfpsclr <= '0';
when s11593 => state := s11594; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (582, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11594 => state := s11595; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1102, 12)); -- offset LSB 1054
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s11595 => state := s11596;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1103, 12)); -- offset MSB 1055
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11596 => state := s11597; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11597 => 			--4
	if (fixed2floatrdy = '1') then state := s11598;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11597; end if;
when s11598 => state := s11599; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11599 => 			--6
	if (mulfprdy = '1') then state := s11600;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11599; end if;
when s11600 => state := s11601; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11601 => 			--8
	if (mulfprdy = '1') then state := s11602;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11601; end if;
when s11602 => state := s11603; 	--9
	mulfpsclr <= '0';
when s11603 => state := s11604; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11604 => 			--11
	if (mulfprdy = '1') then state := s11605;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11604; end if;
when s11605 => state := s11606; 	--12
	mulfpsclr <= '0';
when s11606 => state := s11607; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11607 => 			--14
	if (addfprdy = '1') then state := s11608;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11607; end if;
when s11608 => state := s11609; 	--15
	addfpsclr <= '0';
when s11609 => state := s11610; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11610 => 			--17
	if (addfprdy = '1') then state := s11611;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11610; end if;
when s11611 => state := s11612; 	--18
	addfpsclr <= '0';
when s11612 => state := s11613; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11613 => 			--20
	if (addfprdy = '1') then state := s11614;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11613; end if;
when s11614 => state := s11615; 	--21
	addfpsclr <= '0';
when s11615 => state := s11616; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (583, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11616 => state := s11617; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1104, 12)); -- offset LSB 1056
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s11617 => state := s11618;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1105, 12)); -- offset MSB 1057
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11618 => state := s11619; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11619 => 			--4
	if (fixed2floatrdy = '1') then state := s11620;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11619; end if;
when s11620 => state := s11621; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11621 => 			--6
	if (mulfprdy = '1') then state := s11622;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11621; end if;
when s11622 => state := s11623; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11623 => 			--8
	if (mulfprdy = '1') then state := s11624;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11623; end if;
when s11624 => state := s11625; 	--9
	mulfpsclr <= '0';
when s11625 => state := s11626; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11626 => 			--11
	if (mulfprdy = '1') then state := s11627;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11626; end if;
when s11627 => state := s11628; 	--12
	mulfpsclr <= '0';
when s11628 => state := s11629; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11629 => 			--14
	if (addfprdy = '1') then state := s11630;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11629; end if;
when s11630 => state := s11631; 	--15
	addfpsclr <= '0';
when s11631 => state := s11632; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11632 => 			--17
	if (addfprdy = '1') then state := s11633;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11632; end if;
when s11633 => state := s11634; 	--18
	addfpsclr <= '0';
when s11634 => state := s11635; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11635 => 			--20
	if (addfprdy = '1') then state := s11636;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11635; end if;
when s11636 => state := s11637; 	--21
	addfpsclr <= '0';
when s11637 => state := s11638; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (584, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11638 => state := s11639; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1106, 12)); -- offset LSB 1058
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s11639 => state := s11640;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1107, 12)); -- offset MSB 1059
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11640 => state := s11641; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11641 => 			--4
	if (fixed2floatrdy = '1') then state := s11642;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11641; end if;
when s11642 => state := s11643; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11643 => 			--6
	if (mulfprdy = '1') then state := s11644;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11643; end if;
when s11644 => state := s11645; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11645 => 			--8
	if (mulfprdy = '1') then state := s11646;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11645; end if;
when s11646 => state := s11647; 	--9
	mulfpsclr <= '0';
when s11647 => state := s11648; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11648 => 			--11
	if (mulfprdy = '1') then state := s11649;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11648; end if;
when s11649 => state := s11650; 	--12
	mulfpsclr <= '0';
when s11650 => state := s11651; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11651 => 			--14
	if (addfprdy = '1') then state := s11652;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11651; end if;
when s11652 => state := s11653; 	--15
	addfpsclr <= '0';
when s11653 => state := s11654; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11654 => 			--17
	if (addfprdy = '1') then state := s11655;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11654; end if;
when s11655 => state := s11656; 	--18
	addfpsclr <= '0';
when s11656 => state := s11657; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11657 => 			--20
	if (addfprdy = '1') then state := s11658;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11657; end if;
when s11658 => state := s11659; 	--21
	addfpsclr <= '0';
when s11659 => state := s11660; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (585, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11660 => state := s11661; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1108, 12)); -- offset LSB 1060
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s11661 => state := s11662;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1109, 12)); -- offset MSB 1061
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11662 => state := s11663; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11663 => 			--4
	if (fixed2floatrdy = '1') then state := s11664;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11663; end if;
when s11664 => state := s11665; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11665 => 			--6
	if (mulfprdy = '1') then state := s11666;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11665; end if;
when s11666 => state := s11667; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11667 => 			--8
	if (mulfprdy = '1') then state := s11668;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11667; end if;
when s11668 => state := s11669; 	--9
	mulfpsclr <= '0';
when s11669 => state := s11670; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11670 => 			--11
	if (mulfprdy = '1') then state := s11671;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11670; end if;
when s11671 => state := s11672; 	--12
	mulfpsclr <= '0';
when s11672 => state := s11673; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11673 => 			--14
	if (addfprdy = '1') then state := s11674;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11673; end if;
when s11674 => state := s11675; 	--15
	addfpsclr <= '0';
when s11675 => state := s11676; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11676 => 			--17
	if (addfprdy = '1') then state := s11677;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11676; end if;
when s11677 => state := s11678; 	--18
	addfpsclr <= '0';
when s11678 => state := s11679; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11679 => 			--20
	if (addfprdy = '1') then state := s11680;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11679; end if;
when s11680 => state := s11681; 	--21
	addfpsclr <= '0';
when s11681 => state := s11682; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (586, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11682 => state := s11683; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1110, 12)); -- offset LSB 1062
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s11683 => state := s11684;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1111, 12)); -- offset MSB 1063
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11684 => state := s11685; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11685 => 			--4
	if (fixed2floatrdy = '1') then state := s11686;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11685; end if;
when s11686 => state := s11687; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11687 => 			--6
	if (mulfprdy = '1') then state := s11688;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11687; end if;
when s11688 => state := s11689; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11689 => 			--8
	if (mulfprdy = '1') then state := s11690;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11689; end if;
when s11690 => state := s11691; 	--9
	mulfpsclr <= '0';
when s11691 => state := s11692; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11692 => 			--11
	if (mulfprdy = '1') then state := s11693;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11692; end if;
when s11693 => state := s11694; 	--12
	mulfpsclr <= '0';
when s11694 => state := s11695; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11695 => 			--14
	if (addfprdy = '1') then state := s11696;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11695; end if;
when s11696 => state := s11697; 	--15
	addfpsclr <= '0';
when s11697 => state := s11698; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11698 => 			--17
	if (addfprdy = '1') then state := s11699;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11698; end if;
when s11699 => state := s11700; 	--18
	addfpsclr <= '0';
when s11700 => state := s11701; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11701 => 			--20
	if (addfprdy = '1') then state := s11702;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11701; end if;
when s11702 => state := s11703; 	--21
	addfpsclr <= '0';
when s11703 => state := s11704; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (587, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11704 => state := s11705; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1112, 12)); -- offset LSB 1064
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s11705 => state := s11706;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1113, 12)); -- offset MSB 1065
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11706 => state := s11707; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11707 => 			--4
	if (fixed2floatrdy = '1') then state := s11708;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11707; end if;
when s11708 => state := s11709; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11709 => 			--6
	if (mulfprdy = '1') then state := s11710;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11709; end if;
when s11710 => state := s11711; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11711 => 			--8
	if (mulfprdy = '1') then state := s11712;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11711; end if;
when s11712 => state := s11713; 	--9
	mulfpsclr <= '0';
when s11713 => state := s11714; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11714 => 			--11
	if (mulfprdy = '1') then state := s11715;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11714; end if;
when s11715 => state := s11716; 	--12
	mulfpsclr <= '0';
when s11716 => state := s11717; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11717 => 			--14
	if (addfprdy = '1') then state := s11718;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11717; end if;
when s11718 => state := s11719; 	--15
	addfpsclr <= '0';
when s11719 => state := s11720; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11720 => 			--17
	if (addfprdy = '1') then state := s11721;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11720; end if;
when s11721 => state := s11722; 	--18
	addfpsclr <= '0';
when s11722 => state := s11723; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11723 => 			--20
	if (addfprdy = '1') then state := s11724;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11723; end if;
when s11724 => state := s11725; 	--21
	addfpsclr <= '0';
when s11725 => state := s11726; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (588, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11726 => state := s11727; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1114, 12)); -- offset LSB 1066
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s11727 => state := s11728;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1115, 12)); -- offset MSB 1067
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11728 => state := s11729; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11729 => 			--4
	if (fixed2floatrdy = '1') then state := s11730;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11729; end if;
when s11730 => state := s11731; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11731 => 			--6
	if (mulfprdy = '1') then state := s11732;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11731; end if;
when s11732 => state := s11733; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11733 => 			--8
	if (mulfprdy = '1') then state := s11734;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11733; end if;
when s11734 => state := s11735; 	--9
	mulfpsclr <= '0';
when s11735 => state := s11736; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11736 => 			--11
	if (mulfprdy = '1') then state := s11737;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11736; end if;
when s11737 => state := s11738; 	--12
	mulfpsclr <= '0';
when s11738 => state := s11739; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11739 => 			--14
	if (addfprdy = '1') then state := s11740;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11739; end if;
when s11740 => state := s11741; 	--15
	addfpsclr <= '0';
when s11741 => state := s11742; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11742 => 			--17
	if (addfprdy = '1') then state := s11743;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11742; end if;
when s11743 => state := s11744; 	--18
	addfpsclr <= '0';
when s11744 => state := s11745; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11745 => 			--20
	if (addfprdy = '1') then state := s11746;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11745; end if;
when s11746 => state := s11747; 	--21
	addfpsclr <= '0';
when s11747 => state := s11748; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (589, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11748 => state := s11749; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1116, 12)); -- offset LSB 1068
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s11749 => state := s11750;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1117, 12)); -- offset MSB 1069
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11750 => state := s11751; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11751 => 			--4
	if (fixed2floatrdy = '1') then state := s11752;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11751; end if;
when s11752 => state := s11753; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11753 => 			--6
	if (mulfprdy = '1') then state := s11754;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11753; end if;
when s11754 => state := s11755; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11755 => 			--8
	if (mulfprdy = '1') then state := s11756;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11755; end if;
when s11756 => state := s11757; 	--9
	mulfpsclr <= '0';
when s11757 => state := s11758; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11758 => 			--11
	if (mulfprdy = '1') then state := s11759;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11758; end if;
when s11759 => state := s11760; 	--12
	mulfpsclr <= '0';
when s11760 => state := s11761; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11761 => 			--14
	if (addfprdy = '1') then state := s11762;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11761; end if;
when s11762 => state := s11763; 	--15
	addfpsclr <= '0';
when s11763 => state := s11764; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11764 => 			--17
	if (addfprdy = '1') then state := s11765;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11764; end if;
when s11765 => state := s11766; 	--18
	addfpsclr <= '0';
when s11766 => state := s11767; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11767 => 			--20
	if (addfprdy = '1') then state := s11768;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11767; end if;
when s11768 => state := s11769; 	--21
	addfpsclr <= '0';
when s11769 => state := s11770; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (590, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11770 => state := s11771; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1118, 12)); -- offset LSB 1070
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s11771 => state := s11772;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1119, 12)); -- offset MSB 1071
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11772 => state := s11773; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11773 => 			--4
	if (fixed2floatrdy = '1') then state := s11774;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11773; end if;
when s11774 => state := s11775; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11775 => 			--6
	if (mulfprdy = '1') then state := s11776;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11775; end if;
when s11776 => state := s11777; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11777 => 			--8
	if (mulfprdy = '1') then state := s11778;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11777; end if;
when s11778 => state := s11779; 	--9
	mulfpsclr <= '0';
when s11779 => state := s11780; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11780 => 			--11
	if (mulfprdy = '1') then state := s11781;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11780; end if;
when s11781 => state := s11782; 	--12
	mulfpsclr <= '0';
when s11782 => state := s11783; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11783 => 			--14
	if (addfprdy = '1') then state := s11784;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11783; end if;
when s11784 => state := s11785; 	--15
	addfpsclr <= '0';
when s11785 => state := s11786; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11786 => 			--17
	if (addfprdy = '1') then state := s11787;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11786; end if;
when s11787 => state := s11788; 	--18
	addfpsclr <= '0';
when s11788 => state := s11789; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11789 => 			--20
	if (addfprdy = '1') then state := s11790;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11789; end if;
when s11790 => state := s11791; 	--21
	addfpsclr <= '0';
when s11791 => state := s11792; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (591, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11792 => state := s11793; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1120, 12)); -- offset LSB 1072
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s11793 => state := s11794;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1121, 12)); -- offset MSB 1073
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11794 => state := s11795; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11795 => 			--4
	if (fixed2floatrdy = '1') then state := s11796;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11795; end if;
when s11796 => state := s11797; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11797 => 			--6
	if (mulfprdy = '1') then state := s11798;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11797; end if;
when s11798 => state := s11799; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11799 => 			--8
	if (mulfprdy = '1') then state := s11800;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11799; end if;
when s11800 => state := s11801; 	--9
	mulfpsclr <= '0';
when s11801 => state := s11802; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11802 => 			--11
	if (mulfprdy = '1') then state := s11803;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11802; end if;
when s11803 => state := s11804; 	--12
	mulfpsclr <= '0';
when s11804 => state := s11805; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11805 => 			--14
	if (addfprdy = '1') then state := s11806;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11805; end if;
when s11806 => state := s11807; 	--15
	addfpsclr <= '0';
when s11807 => state := s11808; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11808 => 			--17
	if (addfprdy = '1') then state := s11809;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11808; end if;
when s11809 => state := s11810; 	--18
	addfpsclr <= '0';
when s11810 => state := s11811; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11811 => 			--20
	if (addfprdy = '1') then state := s11812;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11811; end if;
when s11812 => state := s11813; 	--21
	addfpsclr <= '0';
when s11813 => state := s11814; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (592, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11814 => state := s11815; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1122, 12)); -- offset LSB 1074
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s11815 => state := s11816;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1123, 12)); -- offset MSB 1075
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11816 => state := s11817; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11817 => 			--4
	if (fixed2floatrdy = '1') then state := s11818;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11817; end if;
when s11818 => state := s11819; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11819 => 			--6
	if (mulfprdy = '1') then state := s11820;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11819; end if;
when s11820 => state := s11821; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11821 => 			--8
	if (mulfprdy = '1') then state := s11822;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11821; end if;
when s11822 => state := s11823; 	--9
	mulfpsclr <= '0';
when s11823 => state := s11824; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11824 => 			--11
	if (mulfprdy = '1') then state := s11825;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11824; end if;
when s11825 => state := s11826; 	--12
	mulfpsclr <= '0';
when s11826 => state := s11827; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11827 => 			--14
	if (addfprdy = '1') then state := s11828;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11827; end if;
when s11828 => state := s11829; 	--15
	addfpsclr <= '0';
when s11829 => state := s11830; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11830 => 			--17
	if (addfprdy = '1') then state := s11831;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11830; end if;
when s11831 => state := s11832; 	--18
	addfpsclr <= '0';
when s11832 => state := s11833; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11833 => 			--20
	if (addfprdy = '1') then state := s11834;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11833; end if;
when s11834 => state := s11835; 	--21
	addfpsclr <= '0';
when s11835 => state := s11836; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (593, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11836 => state := s11837; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1124, 12)); -- offset LSB 1076
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s11837 => state := s11838;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1125, 12)); -- offset MSB 1077
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11838 => state := s11839; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11839 => 			--4
	if (fixed2floatrdy = '1') then state := s11840;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11839; end if;
when s11840 => state := s11841; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11841 => 			--6
	if (mulfprdy = '1') then state := s11842;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11841; end if;
when s11842 => state := s11843; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11843 => 			--8
	if (mulfprdy = '1') then state := s11844;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11843; end if;
when s11844 => state := s11845; 	--9
	mulfpsclr <= '0';
when s11845 => state := s11846; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11846 => 			--11
	if (mulfprdy = '1') then state := s11847;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11846; end if;
when s11847 => state := s11848; 	--12
	mulfpsclr <= '0';
when s11848 => state := s11849; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11849 => 			--14
	if (addfprdy = '1') then state := s11850;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11849; end if;
when s11850 => state := s11851; 	--15
	addfpsclr <= '0';
when s11851 => state := s11852; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11852 => 			--17
	if (addfprdy = '1') then state := s11853;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11852; end if;
when s11853 => state := s11854; 	--18
	addfpsclr <= '0';
when s11854 => state := s11855; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11855 => 			--20
	if (addfprdy = '1') then state := s11856;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11855; end if;
when s11856 => state := s11857; 	--21
	addfpsclr <= '0';
when s11857 => state := s11858; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (594, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11858 => state := s11859; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1126, 12)); -- offset LSB 1078
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s11859 => state := s11860;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1127, 12)); -- offset MSB 1079
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11860 => state := s11861; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11861 => 			--4
	if (fixed2floatrdy = '1') then state := s11862;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11861; end if;
when s11862 => state := s11863; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11863 => 			--6
	if (mulfprdy = '1') then state := s11864;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11863; end if;
when s11864 => state := s11865; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11865 => 			--8
	if (mulfprdy = '1') then state := s11866;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11865; end if;
when s11866 => state := s11867; 	--9
	mulfpsclr <= '0';
when s11867 => state := s11868; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11868 => 			--11
	if (mulfprdy = '1') then state := s11869;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11868; end if;
when s11869 => state := s11870; 	--12
	mulfpsclr <= '0';
when s11870 => state := s11871; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11871 => 			--14
	if (addfprdy = '1') then state := s11872;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11871; end if;
when s11872 => state := s11873; 	--15
	addfpsclr <= '0';
when s11873 => state := s11874; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11874 => 			--17
	if (addfprdy = '1') then state := s11875;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11874; end if;
when s11875 => state := s11876; 	--18
	addfpsclr <= '0';
when s11876 => state := s11877; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11877 => 			--20
	if (addfprdy = '1') then state := s11878;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11877; end if;
when s11878 => state := s11879; 	--21
	addfpsclr <= '0';
when s11879 => state := s11880; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (595, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11880 => state := s11881; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1128, 12)); -- offset LSB 1080
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s11881 => state := s11882;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1129, 12)); -- offset MSB 1081
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11882 => state := s11883; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11883 => 			--4
	if (fixed2floatrdy = '1') then state := s11884;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11883; end if;
when s11884 => state := s11885; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11885 => 			--6
	if (mulfprdy = '1') then state := s11886;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11885; end if;
when s11886 => state := s11887; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11887 => 			--8
	if (mulfprdy = '1') then state := s11888;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11887; end if;
when s11888 => state := s11889; 	--9
	mulfpsclr <= '0';
when s11889 => state := s11890; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11890 => 			--11
	if (mulfprdy = '1') then state := s11891;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11890; end if;
when s11891 => state := s11892; 	--12
	mulfpsclr <= '0';
when s11892 => state := s11893; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11893 => 			--14
	if (addfprdy = '1') then state := s11894;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11893; end if;
when s11894 => state := s11895; 	--15
	addfpsclr <= '0';
when s11895 => state := s11896; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11896 => 			--17
	if (addfprdy = '1') then state := s11897;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11896; end if;
when s11897 => state := s11898; 	--18
	addfpsclr <= '0';
when s11898 => state := s11899; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11899 => 			--20
	if (addfprdy = '1') then state := s11900;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11899; end if;
when s11900 => state := s11901; 	--21
	addfpsclr <= '0';
when s11901 => state := s11902; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (596, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11902 => state := s11903; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1130, 12)); -- offset LSB 1082
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s11903 => state := s11904;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1131, 12)); -- offset MSB 1083
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11904 => state := s11905; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11905 => 			--4
	if (fixed2floatrdy = '1') then state := s11906;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11905; end if;
when s11906 => state := s11907; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11907 => 			--6
	if (mulfprdy = '1') then state := s11908;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11907; end if;
when s11908 => state := s11909; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11909 => 			--8
	if (mulfprdy = '1') then state := s11910;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11909; end if;
when s11910 => state := s11911; 	--9
	mulfpsclr <= '0';
when s11911 => state := s11912; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11912 => 			--11
	if (mulfprdy = '1') then state := s11913;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11912; end if;
when s11913 => state := s11914; 	--12
	mulfpsclr <= '0';
when s11914 => state := s11915; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11915 => 			--14
	if (addfprdy = '1') then state := s11916;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11915; end if;
when s11916 => state := s11917; 	--15
	addfpsclr <= '0';
when s11917 => state := s11918; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11918 => 			--17
	if (addfprdy = '1') then state := s11919;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11918; end if;
when s11919 => state := s11920; 	--18
	addfpsclr <= '0';
when s11920 => state := s11921; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11921 => 			--20
	if (addfprdy = '1') then state := s11922;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11921; end if;
when s11922 => state := s11923; 	--21
	addfpsclr <= '0';
when s11923 => state := s11924; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (597, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11924 => state := s11925; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1132, 12)); -- offset LSB 1084
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s11925 => state := s11926;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1133, 12)); -- offset MSB 1085
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11926 => state := s11927; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11927 => 			--4
	if (fixed2floatrdy = '1') then state := s11928;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11927; end if;
when s11928 => state := s11929; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11929 => 			--6
	if (mulfprdy = '1') then state := s11930;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11929; end if;
when s11930 => state := s11931; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11931 => 			--8
	if (mulfprdy = '1') then state := s11932;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11931; end if;
when s11932 => state := s11933; 	--9
	mulfpsclr <= '0';
when s11933 => state := s11934; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11934 => 			--11
	if (mulfprdy = '1') then state := s11935;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11934; end if;
when s11935 => state := s11936; 	--12
	mulfpsclr <= '0';
when s11936 => state := s11937; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11937 => 			--14
	if (addfprdy = '1') then state := s11938;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11937; end if;
when s11938 => state := s11939; 	--15
	addfpsclr <= '0';
when s11939 => state := s11940; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11940 => 			--17
	if (addfprdy = '1') then state := s11941;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11940; end if;
when s11941 => state := s11942; 	--18
	addfpsclr <= '0';
when s11942 => state := s11943; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11943 => 			--20
	if (addfprdy = '1') then state := s11944;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11943; end if;
when s11944 => state := s11945; 	--21
	addfpsclr <= '0';
when s11945 => state := s11946; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (598, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11946 => state := s11947; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1134, 12)); -- offset LSB 1086
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s11947 => state := s11948;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1135, 12)); -- offset MSB 1087
	addra <= std_logic_vector (to_unsigned (16, 10)); -- OCCrowI 16
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11948 => state := s11949; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11949 => 			--4
	if (fixed2floatrdy = '1') then state := s11950;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11949; end if;
when s11950 => state := s11951; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11951 => 			--6
	if (mulfprdy = '1') then state := s11952;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11951; end if;
when s11952 => state := s11953; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11953 => 			--8
	if (mulfprdy = '1') then state := s11954;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11953; end if;
when s11954 => state := s11955; 	--9
	mulfpsclr <= '0';
when s11955 => state := s11956; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11956 => 			--11
	if (mulfprdy = '1') then state := s11957;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11956; end if;
when s11957 => state := s11958; 	--12
	mulfpsclr <= '0';
when s11958 => state := s11959; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11959 => 			--14
	if (addfprdy = '1') then state := s11960;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11959; end if;
when s11960 => state := s11961; 	--15
	addfpsclr <= '0';
when s11961 => state := s11962; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11962 => 			--17
	if (addfprdy = '1') then state := s11963;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11962; end if;
when s11963 => state := s11964; 	--18
	addfpsclr <= '0';
when s11964 => state := s11965; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11965 => 			--20
	if (addfprdy = '1') then state := s11966;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11965; end if;
when s11966 => state := s11967; 	--21
	addfpsclr <= '0';
when s11967 => state := s11968; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (599, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11968 => state := s11969; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1136, 12)); -- offset LSB 1088
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s11969 => state := s11970;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1137, 12)); -- offset MSB 1089
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11970 => state := s11971; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11971 => 			--4
	if (fixed2floatrdy = '1') then state := s11972;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11971; end if;
when s11972 => state := s11973; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11973 => 			--6
	if (mulfprdy = '1') then state := s11974;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11973; end if;
when s11974 => state := s11975; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11975 => 			--8
	if (mulfprdy = '1') then state := s11976;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11975; end if;
when s11976 => state := s11977; 	--9
	mulfpsclr <= '0';
when s11977 => state := s11978; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s11978 => 			--11
	if (mulfprdy = '1') then state := s11979;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11978; end if;
when s11979 => state := s11980; 	--12
	mulfpsclr <= '0';
when s11980 => state := s11981; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s11981 => 			--14
	if (addfprdy = '1') then state := s11982;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11981; end if;
when s11982 => state := s11983; 	--15
	addfpsclr <= '0';
when s11983 => state := s11984; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s11984 => 			--17
	if (addfprdy = '1') then state := s11985;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11984; end if;
when s11985 => state := s11986; 	--18
	addfpsclr <= '0';
when s11986 => state := s11987; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s11987 => 			--20
	if (addfprdy = '1') then state := s11988;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s11987; end if;
when s11988 => state := s11989; 	--21
	addfpsclr <= '0';
when s11989 => state := s11990; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (600, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s11990 => state := s11991; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1138, 12)); -- offset LSB 1090
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s11991 => state := s11992;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1139, 12)); -- offset MSB 1091
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s11992 => state := s11993; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s11993 => 			--4
	if (fixed2floatrdy = '1') then state := s11994;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s11993; end if;
when s11994 => state := s11995; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s11995 => 			--6
	if (mulfprdy = '1') then state := s11996;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11995; end if;
when s11996 => state := s11997; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s11997 => 			--8
	if (mulfprdy = '1') then state := s11998;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s11997; end if;
when s11998 => state := s11999; 	--9
	mulfpsclr <= '0';
when s11999 => state := s12000; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12000 => 			--11
	if (mulfprdy = '1') then state := s12001;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12000; end if;
when s12001 => state := s12002; 	--12
	mulfpsclr <= '0';
when s12002 => state := s12003; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12003 => 			--14
	if (addfprdy = '1') then state := s12004;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12003; end if;
when s12004 => state := s12005; 	--15
	addfpsclr <= '0';
when s12005 => state := s12006; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12006 => 			--17
	if (addfprdy = '1') then state := s12007;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12006; end if;
when s12007 => state := s12008; 	--18
	addfpsclr <= '0';
when s12008 => state := s12009; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12009 => 			--20
	if (addfprdy = '1') then state := s12010;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12009; end if;
when s12010 => state := s12011; 	--21
	addfpsclr <= '0';
when s12011 => state := s12012; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (601, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12012 => state := s12013; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1140, 12)); -- offset LSB 1092
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s12013 => state := s12014;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1141, 12)); -- offset MSB 1093
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12014 => state := s12015; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12015 => 			--4
	if (fixed2floatrdy = '1') then state := s12016;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12015; end if;
when s12016 => state := s12017; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12017 => 			--6
	if (mulfprdy = '1') then state := s12018;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12017; end if;
when s12018 => state := s12019; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12019 => 			--8
	if (mulfprdy = '1') then state := s12020;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12019; end if;
when s12020 => state := s12021; 	--9
	mulfpsclr <= '0';
when s12021 => state := s12022; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12022 => 			--11
	if (mulfprdy = '1') then state := s12023;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12022; end if;
when s12023 => state := s12024; 	--12
	mulfpsclr <= '0';
when s12024 => state := s12025; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12025 => 			--14
	if (addfprdy = '1') then state := s12026;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12025; end if;
when s12026 => state := s12027; 	--15
	addfpsclr <= '0';
when s12027 => state := s12028; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12028 => 			--17
	if (addfprdy = '1') then state := s12029;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12028; end if;
when s12029 => state := s12030; 	--18
	addfpsclr <= '0';
when s12030 => state := s12031; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12031 => 			--20
	if (addfprdy = '1') then state := s12032;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12031; end if;
when s12032 => state := s12033; 	--21
	addfpsclr <= '0';
when s12033 => state := s12034; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (602, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12034 => state := s12035; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1142, 12)); -- offset LSB 1094
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s12035 => state := s12036;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1143, 12)); -- offset MSB 1095
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12036 => state := s12037; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12037 => 			--4
	if (fixed2floatrdy = '1') then state := s12038;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12037; end if;
when s12038 => state := s12039; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12039 => 			--6
	if (mulfprdy = '1') then state := s12040;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12039; end if;
when s12040 => state := s12041; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12041 => 			--8
	if (mulfprdy = '1') then state := s12042;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12041; end if;
when s12042 => state := s12043; 	--9
	mulfpsclr <= '0';
when s12043 => state := s12044; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12044 => 			--11
	if (mulfprdy = '1') then state := s12045;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12044; end if;
when s12045 => state := s12046; 	--12
	mulfpsclr <= '0';
when s12046 => state := s12047; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12047 => 			--14
	if (addfprdy = '1') then state := s12048;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12047; end if;
when s12048 => state := s12049; 	--15
	addfpsclr <= '0';
when s12049 => state := s12050; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12050 => 			--17
	if (addfprdy = '1') then state := s12051;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12050; end if;
when s12051 => state := s12052; 	--18
	addfpsclr <= '0';
when s12052 => state := s12053; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12053 => 			--20
	if (addfprdy = '1') then state := s12054;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12053; end if;
when s12054 => state := s12055; 	--21
	addfpsclr <= '0';
when s12055 => state := s12056; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (603, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12056 => state := s12057; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1144, 12)); -- offset LSB 1096
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s12057 => state := s12058;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1145, 12)); -- offset MSB 1097
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12058 => state := s12059; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12059 => 			--4
	if (fixed2floatrdy = '1') then state := s12060;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12059; end if;
when s12060 => state := s12061; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12061 => 			--6
	if (mulfprdy = '1') then state := s12062;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12061; end if;
when s12062 => state := s12063; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12063 => 			--8
	if (mulfprdy = '1') then state := s12064;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12063; end if;
when s12064 => state := s12065; 	--9
	mulfpsclr <= '0';
when s12065 => state := s12066; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12066 => 			--11
	if (mulfprdy = '1') then state := s12067;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12066; end if;
when s12067 => state := s12068; 	--12
	mulfpsclr <= '0';
when s12068 => state := s12069; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12069 => 			--14
	if (addfprdy = '1') then state := s12070;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12069; end if;
when s12070 => state := s12071; 	--15
	addfpsclr <= '0';
when s12071 => state := s12072; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12072 => 			--17
	if (addfprdy = '1') then state := s12073;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12072; end if;
when s12073 => state := s12074; 	--18
	addfpsclr <= '0';
when s12074 => state := s12075; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12075 => 			--20
	if (addfprdy = '1') then state := s12076;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12075; end if;
when s12076 => state := s12077; 	--21
	addfpsclr <= '0';
when s12077 => state := s12078; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (604, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12078 => state := s12079; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1146, 12)); -- offset LSB 1098
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s12079 => state := s12080;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1147, 12)); -- offset MSB 1099
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12080 => state := s12081; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12081 => 			--4
	if (fixed2floatrdy = '1') then state := s12082;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12081; end if;
when s12082 => state := s12083; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12083 => 			--6
	if (mulfprdy = '1') then state := s12084;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12083; end if;
when s12084 => state := s12085; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12085 => 			--8
	if (mulfprdy = '1') then state := s12086;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12085; end if;
when s12086 => state := s12087; 	--9
	mulfpsclr <= '0';
when s12087 => state := s12088; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12088 => 			--11
	if (mulfprdy = '1') then state := s12089;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12088; end if;
when s12089 => state := s12090; 	--12
	mulfpsclr <= '0';
when s12090 => state := s12091; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12091 => 			--14
	if (addfprdy = '1') then state := s12092;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12091; end if;
when s12092 => state := s12093; 	--15
	addfpsclr <= '0';
when s12093 => state := s12094; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12094 => 			--17
	if (addfprdy = '1') then state := s12095;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12094; end if;
when s12095 => state := s12096; 	--18
	addfpsclr <= '0';
when s12096 => state := s12097; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12097 => 			--20
	if (addfprdy = '1') then state := s12098;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12097; end if;
when s12098 => state := s12099; 	--21
	addfpsclr <= '0';
when s12099 => state := s12100; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (605, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12100 => state := s12101; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1148, 12)); -- offset LSB 1100
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s12101 => state := s12102;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1149, 12)); -- offset MSB 1101
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12102 => state := s12103; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12103 => 			--4
	if (fixed2floatrdy = '1') then state := s12104;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12103; end if;
when s12104 => state := s12105; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12105 => 			--6
	if (mulfprdy = '1') then state := s12106;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12105; end if;
when s12106 => state := s12107; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12107 => 			--8
	if (mulfprdy = '1') then state := s12108;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12107; end if;
when s12108 => state := s12109; 	--9
	mulfpsclr <= '0';
when s12109 => state := s12110; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12110 => 			--11
	if (mulfprdy = '1') then state := s12111;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12110; end if;
when s12111 => state := s12112; 	--12
	mulfpsclr <= '0';
when s12112 => state := s12113; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12113 => 			--14
	if (addfprdy = '1') then state := s12114;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12113; end if;
when s12114 => state := s12115; 	--15
	addfpsclr <= '0';
when s12115 => state := s12116; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12116 => 			--17
	if (addfprdy = '1') then state := s12117;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12116; end if;
when s12117 => state := s12118; 	--18
	addfpsclr <= '0';
when s12118 => state := s12119; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12119 => 			--20
	if (addfprdy = '1') then state := s12120;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12119; end if;
when s12120 => state := s12121; 	--21
	addfpsclr <= '0';
when s12121 => state := s12122; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (606, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12122 => state := s12123; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1150, 12)); -- offset LSB 1102
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s12123 => state := s12124;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1151, 12)); -- offset MSB 1103
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12124 => state := s12125; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12125 => 			--4
	if (fixed2floatrdy = '1') then state := s12126;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12125; end if;
when s12126 => state := s12127; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12127 => 			--6
	if (mulfprdy = '1') then state := s12128;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12127; end if;
when s12128 => state := s12129; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12129 => 			--8
	if (mulfprdy = '1') then state := s12130;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12129; end if;
when s12130 => state := s12131; 	--9
	mulfpsclr <= '0';
when s12131 => state := s12132; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12132 => 			--11
	if (mulfprdy = '1') then state := s12133;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12132; end if;
when s12133 => state := s12134; 	--12
	mulfpsclr <= '0';
when s12134 => state := s12135; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12135 => 			--14
	if (addfprdy = '1') then state := s12136;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12135; end if;
when s12136 => state := s12137; 	--15
	addfpsclr <= '0';
when s12137 => state := s12138; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12138 => 			--17
	if (addfprdy = '1') then state := s12139;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12138; end if;
when s12139 => state := s12140; 	--18
	addfpsclr <= '0';
when s12140 => state := s12141; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12141 => 			--20
	if (addfprdy = '1') then state := s12142;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12141; end if;
when s12142 => state := s12143; 	--21
	addfpsclr <= '0';
when s12143 => state := s12144; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (607, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12144 => state := s12145; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1152, 12)); -- offset LSB 1104
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s12145 => state := s12146;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1153, 12)); -- offset MSB 1105
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12146 => state := s12147; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12147 => 			--4
	if (fixed2floatrdy = '1') then state := s12148;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12147; end if;
when s12148 => state := s12149; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12149 => 			--6
	if (mulfprdy = '1') then state := s12150;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12149; end if;
when s12150 => state := s12151; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12151 => 			--8
	if (mulfprdy = '1') then state := s12152;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12151; end if;
when s12152 => state := s12153; 	--9
	mulfpsclr <= '0';
when s12153 => state := s12154; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12154 => 			--11
	if (mulfprdy = '1') then state := s12155;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12154; end if;
when s12155 => state := s12156; 	--12
	mulfpsclr <= '0';
when s12156 => state := s12157; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12157 => 			--14
	if (addfprdy = '1') then state := s12158;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12157; end if;
when s12158 => state := s12159; 	--15
	addfpsclr <= '0';
when s12159 => state := s12160; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12160 => 			--17
	if (addfprdy = '1') then state := s12161;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12160; end if;
when s12161 => state := s12162; 	--18
	addfpsclr <= '0';
when s12162 => state := s12163; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12163 => 			--20
	if (addfprdy = '1') then state := s12164;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12163; end if;
when s12164 => state := s12165; 	--21
	addfpsclr <= '0';
when s12165 => state := s12166; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (608, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12166 => state := s12167; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1154, 12)); -- offset LSB 1106
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s12167 => state := s12168;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1155, 12)); -- offset MSB 1107
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12168 => state := s12169; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12169 => 			--4
	if (fixed2floatrdy = '1') then state := s12170;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12169; end if;
when s12170 => state := s12171; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12171 => 			--6
	if (mulfprdy = '1') then state := s12172;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12171; end if;
when s12172 => state := s12173; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12173 => 			--8
	if (mulfprdy = '1') then state := s12174;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12173; end if;
when s12174 => state := s12175; 	--9
	mulfpsclr <= '0';
when s12175 => state := s12176; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12176 => 			--11
	if (mulfprdy = '1') then state := s12177;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12176; end if;
when s12177 => state := s12178; 	--12
	mulfpsclr <= '0';
when s12178 => state := s12179; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12179 => 			--14
	if (addfprdy = '1') then state := s12180;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12179; end if;
when s12180 => state := s12181; 	--15
	addfpsclr <= '0';
when s12181 => state := s12182; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12182 => 			--17
	if (addfprdy = '1') then state := s12183;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12182; end if;
when s12183 => state := s12184; 	--18
	addfpsclr <= '0';
when s12184 => state := s12185; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12185 => 			--20
	if (addfprdy = '1') then state := s12186;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12185; end if;
when s12186 => state := s12187; 	--21
	addfpsclr <= '0';
when s12187 => state := s12188; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (609, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12188 => state := s12189; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1156, 12)); -- offset LSB 1108
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s12189 => state := s12190;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1157, 12)); -- offset MSB 1109
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12190 => state := s12191; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12191 => 			--4
	if (fixed2floatrdy = '1') then state := s12192;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12191; end if;
when s12192 => state := s12193; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12193 => 			--6
	if (mulfprdy = '1') then state := s12194;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12193; end if;
when s12194 => state := s12195; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12195 => 			--8
	if (mulfprdy = '1') then state := s12196;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12195; end if;
when s12196 => state := s12197; 	--9
	mulfpsclr <= '0';
when s12197 => state := s12198; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12198 => 			--11
	if (mulfprdy = '1') then state := s12199;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12198; end if;
when s12199 => state := s12200; 	--12
	mulfpsclr <= '0';
when s12200 => state := s12201; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12201 => 			--14
	if (addfprdy = '1') then state := s12202;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12201; end if;
when s12202 => state := s12203; 	--15
	addfpsclr <= '0';
when s12203 => state := s12204; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12204 => 			--17
	if (addfprdy = '1') then state := s12205;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12204; end if;
when s12205 => state := s12206; 	--18
	addfpsclr <= '0';
when s12206 => state := s12207; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12207 => 			--20
	if (addfprdy = '1') then state := s12208;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12207; end if;
when s12208 => state := s12209; 	--21
	addfpsclr <= '0';
when s12209 => state := s12210; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (610, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12210 => state := s12211; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1158, 12)); -- offset LSB 1110
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s12211 => state := s12212;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1159, 12)); -- offset MSB 1111
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12212 => state := s12213; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12213 => 			--4
	if (fixed2floatrdy = '1') then state := s12214;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12213; end if;
when s12214 => state := s12215; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12215 => 			--6
	if (mulfprdy = '1') then state := s12216;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12215; end if;
when s12216 => state := s12217; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12217 => 			--8
	if (mulfprdy = '1') then state := s12218;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12217; end if;
when s12218 => state := s12219; 	--9
	mulfpsclr <= '0';
when s12219 => state := s12220; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12220 => 			--11
	if (mulfprdy = '1') then state := s12221;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12220; end if;
when s12221 => state := s12222; 	--12
	mulfpsclr <= '0';
when s12222 => state := s12223; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12223 => 			--14
	if (addfprdy = '1') then state := s12224;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12223; end if;
when s12224 => state := s12225; 	--15
	addfpsclr <= '0';
when s12225 => state := s12226; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12226 => 			--17
	if (addfprdy = '1') then state := s12227;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12226; end if;
when s12227 => state := s12228; 	--18
	addfpsclr <= '0';
when s12228 => state := s12229; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12229 => 			--20
	if (addfprdy = '1') then state := s12230;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12229; end if;
when s12230 => state := s12231; 	--21
	addfpsclr <= '0';
when s12231 => state := s12232; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (611, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12232 => state := s12233; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1160, 12)); -- offset LSB 1112
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s12233 => state := s12234;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1161, 12)); -- offset MSB 1113
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12234 => state := s12235; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12235 => 			--4
	if (fixed2floatrdy = '1') then state := s12236;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12235; end if;
when s12236 => state := s12237; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12237 => 			--6
	if (mulfprdy = '1') then state := s12238;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12237; end if;
when s12238 => state := s12239; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12239 => 			--8
	if (mulfprdy = '1') then state := s12240;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12239; end if;
when s12240 => state := s12241; 	--9
	mulfpsclr <= '0';
when s12241 => state := s12242; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12242 => 			--11
	if (mulfprdy = '1') then state := s12243;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12242; end if;
when s12243 => state := s12244; 	--12
	mulfpsclr <= '0';
when s12244 => state := s12245; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12245 => 			--14
	if (addfprdy = '1') then state := s12246;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12245; end if;
when s12246 => state := s12247; 	--15
	addfpsclr <= '0';
when s12247 => state := s12248; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12248 => 			--17
	if (addfprdy = '1') then state := s12249;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12248; end if;
when s12249 => state := s12250; 	--18
	addfpsclr <= '0';
when s12250 => state := s12251; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12251 => 			--20
	if (addfprdy = '1') then state := s12252;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12251; end if;
when s12252 => state := s12253; 	--21
	addfpsclr <= '0';
when s12253 => state := s12254; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (612, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12254 => state := s12255; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1162, 12)); -- offset LSB 1114
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s12255 => state := s12256;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1163, 12)); -- offset MSB 1115
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12256 => state := s12257; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12257 => 			--4
	if (fixed2floatrdy = '1') then state := s12258;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12257; end if;
when s12258 => state := s12259; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12259 => 			--6
	if (mulfprdy = '1') then state := s12260;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12259; end if;
when s12260 => state := s12261; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12261 => 			--8
	if (mulfprdy = '1') then state := s12262;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12261; end if;
when s12262 => state := s12263; 	--9
	mulfpsclr <= '0';
when s12263 => state := s12264; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12264 => 			--11
	if (mulfprdy = '1') then state := s12265;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12264; end if;
when s12265 => state := s12266; 	--12
	mulfpsclr <= '0';
when s12266 => state := s12267; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12267 => 			--14
	if (addfprdy = '1') then state := s12268;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12267; end if;
when s12268 => state := s12269; 	--15
	addfpsclr <= '0';
when s12269 => state := s12270; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12270 => 			--17
	if (addfprdy = '1') then state := s12271;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12270; end if;
when s12271 => state := s12272; 	--18
	addfpsclr <= '0';
when s12272 => state := s12273; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12273 => 			--20
	if (addfprdy = '1') then state := s12274;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12273; end if;
when s12274 => state := s12275; 	--21
	addfpsclr <= '0';
when s12275 => state := s12276; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (613, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12276 => state := s12277; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1164, 12)); -- offset LSB 1116
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s12277 => state := s12278;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1165, 12)); -- offset MSB 1117
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12278 => state := s12279; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12279 => 			--4
	if (fixed2floatrdy = '1') then state := s12280;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12279; end if;
when s12280 => state := s12281; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12281 => 			--6
	if (mulfprdy = '1') then state := s12282;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12281; end if;
when s12282 => state := s12283; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12283 => 			--8
	if (mulfprdy = '1') then state := s12284;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12283; end if;
when s12284 => state := s12285; 	--9
	mulfpsclr <= '0';
when s12285 => state := s12286; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12286 => 			--11
	if (mulfprdy = '1') then state := s12287;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12286; end if;
when s12287 => state := s12288; 	--12
	mulfpsclr <= '0';
when s12288 => state := s12289; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12289 => 			--14
	if (addfprdy = '1') then state := s12290;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12289; end if;
when s12290 => state := s12291; 	--15
	addfpsclr <= '0';
when s12291 => state := s12292; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12292 => 			--17
	if (addfprdy = '1') then state := s12293;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12292; end if;
when s12293 => state := s12294; 	--18
	addfpsclr <= '0';
when s12294 => state := s12295; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12295 => 			--20
	if (addfprdy = '1') then state := s12296;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12295; end if;
when s12296 => state := s12297; 	--21
	addfpsclr <= '0';
when s12297 => state := s12298; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (614, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12298 => state := s12299; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1166, 12)); -- offset LSB 1118
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s12299 => state := s12300;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1167, 12)); -- offset MSB 1119
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12300 => state := s12301; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12301 => 			--4
	if (fixed2floatrdy = '1') then state := s12302;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12301; end if;
when s12302 => state := s12303; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12303 => 			--6
	if (mulfprdy = '1') then state := s12304;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12303; end if;
when s12304 => state := s12305; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12305 => 			--8
	if (mulfprdy = '1') then state := s12306;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12305; end if;
when s12306 => state := s12307; 	--9
	mulfpsclr <= '0';
when s12307 => state := s12308; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12308 => 			--11
	if (mulfprdy = '1') then state := s12309;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12308; end if;
when s12309 => state := s12310; 	--12
	mulfpsclr <= '0';
when s12310 => state := s12311; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12311 => 			--14
	if (addfprdy = '1') then state := s12312;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12311; end if;
when s12312 => state := s12313; 	--15
	addfpsclr <= '0';
when s12313 => state := s12314; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12314 => 			--17
	if (addfprdy = '1') then state := s12315;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12314; end if;
when s12315 => state := s12316; 	--18
	addfpsclr <= '0';
when s12316 => state := s12317; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12317 => 			--20
	if (addfprdy = '1') then state := s12318;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12317; end if;
when s12318 => state := s12319; 	--21
	addfpsclr <= '0';
when s12319 => state := s12320; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (615, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12320 => state := s12321; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1168, 12)); -- offset LSB 1120
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s12321 => state := s12322;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1169, 12)); -- offset MSB 1121
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12322 => state := s12323; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12323 => 			--4
	if (fixed2floatrdy = '1') then state := s12324;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12323; end if;
when s12324 => state := s12325; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12325 => 			--6
	if (mulfprdy = '1') then state := s12326;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12325; end if;
when s12326 => state := s12327; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12327 => 			--8
	if (mulfprdy = '1') then state := s12328;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12327; end if;
when s12328 => state := s12329; 	--9
	mulfpsclr <= '0';
when s12329 => state := s12330; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12330 => 			--11
	if (mulfprdy = '1') then state := s12331;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12330; end if;
when s12331 => state := s12332; 	--12
	mulfpsclr <= '0';
when s12332 => state := s12333; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12333 => 			--14
	if (addfprdy = '1') then state := s12334;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12333; end if;
when s12334 => state := s12335; 	--15
	addfpsclr <= '0';
when s12335 => state := s12336; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12336 => 			--17
	if (addfprdy = '1') then state := s12337;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12336; end if;
when s12337 => state := s12338; 	--18
	addfpsclr <= '0';
when s12338 => state := s12339; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12339 => 			--20
	if (addfprdy = '1') then state := s12340;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12339; end if;
when s12340 => state := s12341; 	--21
	addfpsclr <= '0';
when s12341 => state := s12342; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (616, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12342 => state := s12343; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1170, 12)); -- offset LSB 1122
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s12343 => state := s12344;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1171, 12)); -- offset MSB 1123
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12344 => state := s12345; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12345 => 			--4
	if (fixed2floatrdy = '1') then state := s12346;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12345; end if;
when s12346 => state := s12347; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12347 => 			--6
	if (mulfprdy = '1') then state := s12348;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12347; end if;
when s12348 => state := s12349; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12349 => 			--8
	if (mulfprdy = '1') then state := s12350;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12349; end if;
when s12350 => state := s12351; 	--9
	mulfpsclr <= '0';
when s12351 => state := s12352; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12352 => 			--11
	if (mulfprdy = '1') then state := s12353;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12352; end if;
when s12353 => state := s12354; 	--12
	mulfpsclr <= '0';
when s12354 => state := s12355; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12355 => 			--14
	if (addfprdy = '1') then state := s12356;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12355; end if;
when s12356 => state := s12357; 	--15
	addfpsclr <= '0';
when s12357 => state := s12358; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12358 => 			--17
	if (addfprdy = '1') then state := s12359;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12358; end if;
when s12359 => state := s12360; 	--18
	addfpsclr <= '0';
when s12360 => state := s12361; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12361 => 			--20
	if (addfprdy = '1') then state := s12362;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12361; end if;
when s12362 => state := s12363; 	--21
	addfpsclr <= '0';
when s12363 => state := s12364; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (617, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12364 => state := s12365; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1172, 12)); -- offset LSB 1124
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s12365 => state := s12366;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1173, 12)); -- offset MSB 1125
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12366 => state := s12367; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12367 => 			--4
	if (fixed2floatrdy = '1') then state := s12368;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12367; end if;
when s12368 => state := s12369; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12369 => 			--6
	if (mulfprdy = '1') then state := s12370;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12369; end if;
when s12370 => state := s12371; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12371 => 			--8
	if (mulfprdy = '1') then state := s12372;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12371; end if;
when s12372 => state := s12373; 	--9
	mulfpsclr <= '0';
when s12373 => state := s12374; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12374 => 			--11
	if (mulfprdy = '1') then state := s12375;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12374; end if;
when s12375 => state := s12376; 	--12
	mulfpsclr <= '0';
when s12376 => state := s12377; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12377 => 			--14
	if (addfprdy = '1') then state := s12378;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12377; end if;
when s12378 => state := s12379; 	--15
	addfpsclr <= '0';
when s12379 => state := s12380; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12380 => 			--17
	if (addfprdy = '1') then state := s12381;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12380; end if;
when s12381 => state := s12382; 	--18
	addfpsclr <= '0';
when s12382 => state := s12383; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12383 => 			--20
	if (addfprdy = '1') then state := s12384;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12383; end if;
when s12384 => state := s12385; 	--21
	addfpsclr <= '0';
when s12385 => state := s12386; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (618, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12386 => state := s12387; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1174, 12)); -- offset LSB 1126
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s12387 => state := s12388;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1175, 12)); -- offset MSB 1127
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12388 => state := s12389; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12389 => 			--4
	if (fixed2floatrdy = '1') then state := s12390;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12389; end if;
when s12390 => state := s12391; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12391 => 			--6
	if (mulfprdy = '1') then state := s12392;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12391; end if;
when s12392 => state := s12393; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12393 => 			--8
	if (mulfprdy = '1') then state := s12394;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12393; end if;
when s12394 => state := s12395; 	--9
	mulfpsclr <= '0';
when s12395 => state := s12396; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12396 => 			--11
	if (mulfprdy = '1') then state := s12397;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12396; end if;
when s12397 => state := s12398; 	--12
	mulfpsclr <= '0';
when s12398 => state := s12399; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12399 => 			--14
	if (addfprdy = '1') then state := s12400;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12399; end if;
when s12400 => state := s12401; 	--15
	addfpsclr <= '0';
when s12401 => state := s12402; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12402 => 			--17
	if (addfprdy = '1') then state := s12403;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12402; end if;
when s12403 => state := s12404; 	--18
	addfpsclr <= '0';
when s12404 => state := s12405; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12405 => 			--20
	if (addfprdy = '1') then state := s12406;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12405; end if;
when s12406 => state := s12407; 	--21
	addfpsclr <= '0';
when s12407 => state := s12408; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (619, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12408 => state := s12409; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1176, 12)); -- offset LSB 1128
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s12409 => state := s12410;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1177, 12)); -- offset MSB 1129
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12410 => state := s12411; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12411 => 			--4
	if (fixed2floatrdy = '1') then state := s12412;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12411; end if;
when s12412 => state := s12413; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12413 => 			--6
	if (mulfprdy = '1') then state := s12414;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12413; end if;
when s12414 => state := s12415; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12415 => 			--8
	if (mulfprdy = '1') then state := s12416;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12415; end if;
when s12416 => state := s12417; 	--9
	mulfpsclr <= '0';
when s12417 => state := s12418; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12418 => 			--11
	if (mulfprdy = '1') then state := s12419;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12418; end if;
when s12419 => state := s12420; 	--12
	mulfpsclr <= '0';
when s12420 => state := s12421; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12421 => 			--14
	if (addfprdy = '1') then state := s12422;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12421; end if;
when s12422 => state := s12423; 	--15
	addfpsclr <= '0';
when s12423 => state := s12424; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12424 => 			--17
	if (addfprdy = '1') then state := s12425;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12424; end if;
when s12425 => state := s12426; 	--18
	addfpsclr <= '0';
when s12426 => state := s12427; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12427 => 			--20
	if (addfprdy = '1') then state := s12428;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12427; end if;
when s12428 => state := s12429; 	--21
	addfpsclr <= '0';
when s12429 => state := s12430; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (620, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12430 => state := s12431; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1178, 12)); -- offset LSB 1130
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s12431 => state := s12432;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1179, 12)); -- offset MSB 1131
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12432 => state := s12433; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12433 => 			--4
	if (fixed2floatrdy = '1') then state := s12434;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12433; end if;
when s12434 => state := s12435; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12435 => 			--6
	if (mulfprdy = '1') then state := s12436;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12435; end if;
when s12436 => state := s12437; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12437 => 			--8
	if (mulfprdy = '1') then state := s12438;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12437; end if;
when s12438 => state := s12439; 	--9
	mulfpsclr <= '0';
when s12439 => state := s12440; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12440 => 			--11
	if (mulfprdy = '1') then state := s12441;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12440; end if;
when s12441 => state := s12442; 	--12
	mulfpsclr <= '0';
when s12442 => state := s12443; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12443 => 			--14
	if (addfprdy = '1') then state := s12444;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12443; end if;
when s12444 => state := s12445; 	--15
	addfpsclr <= '0';
when s12445 => state := s12446; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12446 => 			--17
	if (addfprdy = '1') then state := s12447;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12446; end if;
when s12447 => state := s12448; 	--18
	addfpsclr <= '0';
when s12448 => state := s12449; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12449 => 			--20
	if (addfprdy = '1') then state := s12450;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12449; end if;
when s12450 => state := s12451; 	--21
	addfpsclr <= '0';
when s12451 => state := s12452; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (621, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12452 => state := s12453; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1180, 12)); -- offset LSB 1132
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s12453 => state := s12454;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1181, 12)); -- offset MSB 1133
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12454 => state := s12455; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12455 => 			--4
	if (fixed2floatrdy = '1') then state := s12456;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12455; end if;
when s12456 => state := s12457; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12457 => 			--6
	if (mulfprdy = '1') then state := s12458;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12457; end if;
when s12458 => state := s12459; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12459 => 			--8
	if (mulfprdy = '1') then state := s12460;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12459; end if;
when s12460 => state := s12461; 	--9
	mulfpsclr <= '0';
when s12461 => state := s12462; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12462 => 			--11
	if (mulfprdy = '1') then state := s12463;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12462; end if;
when s12463 => state := s12464; 	--12
	mulfpsclr <= '0';
when s12464 => state := s12465; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12465 => 			--14
	if (addfprdy = '1') then state := s12466;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12465; end if;
when s12466 => state := s12467; 	--15
	addfpsclr <= '0';
when s12467 => state := s12468; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12468 => 			--17
	if (addfprdy = '1') then state := s12469;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12468; end if;
when s12469 => state := s12470; 	--18
	addfpsclr <= '0';
when s12470 => state := s12471; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12471 => 			--20
	if (addfprdy = '1') then state := s12472;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12471; end if;
when s12472 => state := s12473; 	--21
	addfpsclr <= '0';
when s12473 => state := s12474; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (622, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12474 => state := s12475; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1182, 12)); -- offset LSB 1134
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s12475 => state := s12476;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1183, 12)); -- offset MSB 1135
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12476 => state := s12477; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12477 => 			--4
	if (fixed2floatrdy = '1') then state := s12478;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12477; end if;
when s12478 => state := s12479; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12479 => 			--6
	if (mulfprdy = '1') then state := s12480;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12479; end if;
when s12480 => state := s12481; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12481 => 			--8
	if (mulfprdy = '1') then state := s12482;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12481; end if;
when s12482 => state := s12483; 	--9
	mulfpsclr <= '0';
when s12483 => state := s12484; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12484 => 			--11
	if (mulfprdy = '1') then state := s12485;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12484; end if;
when s12485 => state := s12486; 	--12
	mulfpsclr <= '0';
when s12486 => state := s12487; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12487 => 			--14
	if (addfprdy = '1') then state := s12488;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12487; end if;
when s12488 => state := s12489; 	--15
	addfpsclr <= '0';
when s12489 => state := s12490; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12490 => 			--17
	if (addfprdy = '1') then state := s12491;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12490; end if;
when s12491 => state := s12492; 	--18
	addfpsclr <= '0';
when s12492 => state := s12493; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12493 => 			--20
	if (addfprdy = '1') then state := s12494;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12493; end if;
when s12494 => state := s12495; 	--21
	addfpsclr <= '0';
when s12495 => state := s12496; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (623, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12496 => state := s12497; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1184, 12)); -- offset LSB 1136
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s12497 => state := s12498;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1185, 12)); -- offset MSB 1137
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12498 => state := s12499; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12499 => 			--4
	if (fixed2floatrdy = '1') then state := s12500;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12499; end if;
when s12500 => state := s12501; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12501 => 			--6
	if (mulfprdy = '1') then state := s12502;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12501; end if;
when s12502 => state := s12503; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12503 => 			--8
	if (mulfprdy = '1') then state := s12504;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12503; end if;
when s12504 => state := s12505; 	--9
	mulfpsclr <= '0';
when s12505 => state := s12506; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12506 => 			--11
	if (mulfprdy = '1') then state := s12507;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12506; end if;
when s12507 => state := s12508; 	--12
	mulfpsclr <= '0';
when s12508 => state := s12509; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12509 => 			--14
	if (addfprdy = '1') then state := s12510;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12509; end if;
when s12510 => state := s12511; 	--15
	addfpsclr <= '0';
when s12511 => state := s12512; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12512 => 			--17
	if (addfprdy = '1') then state := s12513;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12512; end if;
when s12513 => state := s12514; 	--18
	addfpsclr <= '0';
when s12514 => state := s12515; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12515 => 			--20
	if (addfprdy = '1') then state := s12516;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12515; end if;
when s12516 => state := s12517; 	--21
	addfpsclr <= '0';
when s12517 => state := s12518; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (624, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12518 => state := s12519; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1186, 12)); -- offset LSB 1138
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s12519 => state := s12520;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1187, 12)); -- offset MSB 1139
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12520 => state := s12521; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12521 => 			--4
	if (fixed2floatrdy = '1') then state := s12522;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12521; end if;
when s12522 => state := s12523; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12523 => 			--6
	if (mulfprdy = '1') then state := s12524;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12523; end if;
when s12524 => state := s12525; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12525 => 			--8
	if (mulfprdy = '1') then state := s12526;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12525; end if;
when s12526 => state := s12527; 	--9
	mulfpsclr <= '0';
when s12527 => state := s12528; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12528 => 			--11
	if (mulfprdy = '1') then state := s12529;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12528; end if;
when s12529 => state := s12530; 	--12
	mulfpsclr <= '0';
when s12530 => state := s12531; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12531 => 			--14
	if (addfprdy = '1') then state := s12532;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12531; end if;
when s12532 => state := s12533; 	--15
	addfpsclr <= '0';
when s12533 => state := s12534; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12534 => 			--17
	if (addfprdy = '1') then state := s12535;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12534; end if;
when s12535 => state := s12536; 	--18
	addfpsclr <= '0';
when s12536 => state := s12537; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12537 => 			--20
	if (addfprdy = '1') then state := s12538;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12537; end if;
when s12538 => state := s12539; 	--21
	addfpsclr <= '0';
when s12539 => state := s12540; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (625, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12540 => state := s12541; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1188, 12)); -- offset LSB 1140
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s12541 => state := s12542;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1189, 12)); -- offset MSB 1141
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12542 => state := s12543; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12543 => 			--4
	if (fixed2floatrdy = '1') then state := s12544;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12543; end if;
when s12544 => state := s12545; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12545 => 			--6
	if (mulfprdy = '1') then state := s12546;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12545; end if;
when s12546 => state := s12547; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12547 => 			--8
	if (mulfprdy = '1') then state := s12548;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12547; end if;
when s12548 => state := s12549; 	--9
	mulfpsclr <= '0';
when s12549 => state := s12550; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12550 => 			--11
	if (mulfprdy = '1') then state := s12551;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12550; end if;
when s12551 => state := s12552; 	--12
	mulfpsclr <= '0';
when s12552 => state := s12553; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12553 => 			--14
	if (addfprdy = '1') then state := s12554;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12553; end if;
when s12554 => state := s12555; 	--15
	addfpsclr <= '0';
when s12555 => state := s12556; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12556 => 			--17
	if (addfprdy = '1') then state := s12557;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12556; end if;
when s12557 => state := s12558; 	--18
	addfpsclr <= '0';
when s12558 => state := s12559; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12559 => 			--20
	if (addfprdy = '1') then state := s12560;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12559; end if;
when s12560 => state := s12561; 	--21
	addfpsclr <= '0';
when s12561 => state := s12562; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (626, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12562 => state := s12563; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1190, 12)); -- offset LSB 1142
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s12563 => state := s12564;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1191, 12)); -- offset MSB 1143
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12564 => state := s12565; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12565 => 			--4
	if (fixed2floatrdy = '1') then state := s12566;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12565; end if;
when s12566 => state := s12567; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12567 => 			--6
	if (mulfprdy = '1') then state := s12568;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12567; end if;
when s12568 => state := s12569; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12569 => 			--8
	if (mulfprdy = '1') then state := s12570;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12569; end if;
when s12570 => state := s12571; 	--9
	mulfpsclr <= '0';
when s12571 => state := s12572; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12572 => 			--11
	if (mulfprdy = '1') then state := s12573;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12572; end if;
when s12573 => state := s12574; 	--12
	mulfpsclr <= '0';
when s12574 => state := s12575; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12575 => 			--14
	if (addfprdy = '1') then state := s12576;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12575; end if;
when s12576 => state := s12577; 	--15
	addfpsclr <= '0';
when s12577 => state := s12578; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12578 => 			--17
	if (addfprdy = '1') then state := s12579;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12578; end if;
when s12579 => state := s12580; 	--18
	addfpsclr <= '0';
when s12580 => state := s12581; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12581 => 			--20
	if (addfprdy = '1') then state := s12582;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12581; end if;
when s12582 => state := s12583; 	--21
	addfpsclr <= '0';
when s12583 => state := s12584; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (627, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12584 => state := s12585; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1192, 12)); -- offset LSB 1144
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s12585 => state := s12586;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1193, 12)); -- offset MSB 1145
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12586 => state := s12587; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12587 => 			--4
	if (fixed2floatrdy = '1') then state := s12588;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12587; end if;
when s12588 => state := s12589; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12589 => 			--6
	if (mulfprdy = '1') then state := s12590;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12589; end if;
when s12590 => state := s12591; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12591 => 			--8
	if (mulfprdy = '1') then state := s12592;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12591; end if;
when s12592 => state := s12593; 	--9
	mulfpsclr <= '0';
when s12593 => state := s12594; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12594 => 			--11
	if (mulfprdy = '1') then state := s12595;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12594; end if;
when s12595 => state := s12596; 	--12
	mulfpsclr <= '0';
when s12596 => state := s12597; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12597 => 			--14
	if (addfprdy = '1') then state := s12598;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12597; end if;
when s12598 => state := s12599; 	--15
	addfpsclr <= '0';
when s12599 => state := s12600; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12600 => 			--17
	if (addfprdy = '1') then state := s12601;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12600; end if;
when s12601 => state := s12602; 	--18
	addfpsclr <= '0';
when s12602 => state := s12603; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12603 => 			--20
	if (addfprdy = '1') then state := s12604;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12603; end if;
when s12604 => state := s12605; 	--21
	addfpsclr <= '0';
when s12605 => state := s12606; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (628, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12606 => state := s12607; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1194, 12)); -- offset LSB 1146
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s12607 => state := s12608;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1195, 12)); -- offset MSB 1147
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12608 => state := s12609; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12609 => 			--4
	if (fixed2floatrdy = '1') then state := s12610;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12609; end if;
when s12610 => state := s12611; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12611 => 			--6
	if (mulfprdy = '1') then state := s12612;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12611; end if;
when s12612 => state := s12613; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12613 => 			--8
	if (mulfprdy = '1') then state := s12614;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12613; end if;
when s12614 => state := s12615; 	--9
	mulfpsclr <= '0';
when s12615 => state := s12616; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12616 => 			--11
	if (mulfprdy = '1') then state := s12617;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12616; end if;
when s12617 => state := s12618; 	--12
	mulfpsclr <= '0';
when s12618 => state := s12619; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12619 => 			--14
	if (addfprdy = '1') then state := s12620;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12619; end if;
when s12620 => state := s12621; 	--15
	addfpsclr <= '0';
when s12621 => state := s12622; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12622 => 			--17
	if (addfprdy = '1') then state := s12623;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12622; end if;
when s12623 => state := s12624; 	--18
	addfpsclr <= '0';
when s12624 => state := s12625; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12625 => 			--20
	if (addfprdy = '1') then state := s12626;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12625; end if;
when s12626 => state := s12627; 	--21
	addfpsclr <= '0';
when s12627 => state := s12628; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (629, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12628 => state := s12629; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1196, 12)); -- offset LSB 1148
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s12629 => state := s12630;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1197, 12)); -- offset MSB 1149
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12630 => state := s12631; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12631 => 			--4
	if (fixed2floatrdy = '1') then state := s12632;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12631; end if;
when s12632 => state := s12633; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12633 => 			--6
	if (mulfprdy = '1') then state := s12634;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12633; end if;
when s12634 => state := s12635; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12635 => 			--8
	if (mulfprdy = '1') then state := s12636;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12635; end if;
when s12636 => state := s12637; 	--9
	mulfpsclr <= '0';
when s12637 => state := s12638; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12638 => 			--11
	if (mulfprdy = '1') then state := s12639;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12638; end if;
when s12639 => state := s12640; 	--12
	mulfpsclr <= '0';
when s12640 => state := s12641; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12641 => 			--14
	if (addfprdy = '1') then state := s12642;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12641; end if;
when s12642 => state := s12643; 	--15
	addfpsclr <= '0';
when s12643 => state := s12644; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12644 => 			--17
	if (addfprdy = '1') then state := s12645;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12644; end if;
when s12645 => state := s12646; 	--18
	addfpsclr <= '0';
when s12646 => state := s12647; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12647 => 			--20
	if (addfprdy = '1') then state := s12648;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12647; end if;
when s12648 => state := s12649; 	--21
	addfpsclr <= '0';
when s12649 => state := s12650; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (630, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12650 => state := s12651; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1198, 12)); -- offset LSB 1150
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s12651 => state := s12652;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1199, 12)); -- offset MSB 1151
	addra <= std_logic_vector (to_unsigned (17, 10)); -- OCCrowI 17
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12652 => state := s12653; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12653 => 			--4
	if (fixed2floatrdy = '1') then state := s12654;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12653; end if;
when s12654 => state := s12655; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12655 => 			--6
	if (mulfprdy = '1') then state := s12656;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12655; end if;
when s12656 => state := s12657; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12657 => 			--8
	if (mulfprdy = '1') then state := s12658;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12657; end if;
when s12658 => state := s12659; 	--9
	mulfpsclr <= '0';
when s12659 => state := s12660; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12660 => 			--11
	if (mulfprdy = '1') then state := s12661;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12660; end if;
when s12661 => state := s12662; 	--12
	mulfpsclr <= '0';
when s12662 => state := s12663; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12663 => 			--14
	if (addfprdy = '1') then state := s12664;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12663; end if;
when s12664 => state := s12665; 	--15
	addfpsclr <= '0';
when s12665 => state := s12666; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12666 => 			--17
	if (addfprdy = '1') then state := s12667;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12666; end if;
when s12667 => state := s12668; 	--18
	addfpsclr <= '0';
when s12668 => state := s12669; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12669 => 			--20
	if (addfprdy = '1') then state := s12670;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12669; end if;
when s12670 => state := s12671; 	--21
	addfpsclr <= '0';
when s12671 => state := s12672; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (631, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12672 => state := s12673; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1200, 12)); -- offset LSB 1152
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s12673 => state := s12674;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1201, 12)); -- offset MSB 1153
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12674 => state := s12675; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12675 => 			--4
	if (fixed2floatrdy = '1') then state := s12676;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12675; end if;
when s12676 => state := s12677; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12677 => 			--6
	if (mulfprdy = '1') then state := s12678;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12677; end if;
when s12678 => state := s12679; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12679 => 			--8
	if (mulfprdy = '1') then state := s12680;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12679; end if;
when s12680 => state := s12681; 	--9
	mulfpsclr <= '0';
when s12681 => state := s12682; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12682 => 			--11
	if (mulfprdy = '1') then state := s12683;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12682; end if;
when s12683 => state := s12684; 	--12
	mulfpsclr <= '0';
when s12684 => state := s12685; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12685 => 			--14
	if (addfprdy = '1') then state := s12686;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12685; end if;
when s12686 => state := s12687; 	--15
	addfpsclr <= '0';
when s12687 => state := s12688; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12688 => 			--17
	if (addfprdy = '1') then state := s12689;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12688; end if;
when s12689 => state := s12690; 	--18
	addfpsclr <= '0';
when s12690 => state := s12691; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12691 => 			--20
	if (addfprdy = '1') then state := s12692;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12691; end if;
when s12692 => state := s12693; 	--21
	addfpsclr <= '0';
when s12693 => state := s12694; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (632, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12694 => state := s12695; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1202, 12)); -- offset LSB 1154
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s12695 => state := s12696;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1203, 12)); -- offset MSB 1155
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12696 => state := s12697; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12697 => 			--4
	if (fixed2floatrdy = '1') then state := s12698;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12697; end if;
when s12698 => state := s12699; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12699 => 			--6
	if (mulfprdy = '1') then state := s12700;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12699; end if;
when s12700 => state := s12701; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12701 => 			--8
	if (mulfprdy = '1') then state := s12702;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12701; end if;
when s12702 => state := s12703; 	--9
	mulfpsclr <= '0';
when s12703 => state := s12704; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12704 => 			--11
	if (mulfprdy = '1') then state := s12705;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12704; end if;
when s12705 => state := s12706; 	--12
	mulfpsclr <= '0';
when s12706 => state := s12707; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12707 => 			--14
	if (addfprdy = '1') then state := s12708;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12707; end if;
when s12708 => state := s12709; 	--15
	addfpsclr <= '0';
when s12709 => state := s12710; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12710 => 			--17
	if (addfprdy = '1') then state := s12711;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12710; end if;
when s12711 => state := s12712; 	--18
	addfpsclr <= '0';
when s12712 => state := s12713; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12713 => 			--20
	if (addfprdy = '1') then state := s12714;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12713; end if;
when s12714 => state := s12715; 	--21
	addfpsclr <= '0';
when s12715 => state := s12716; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (633, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12716 => state := s12717; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1204, 12)); -- offset LSB 1156
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s12717 => state := s12718;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1205, 12)); -- offset MSB 1157
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12718 => state := s12719; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12719 => 			--4
	if (fixed2floatrdy = '1') then state := s12720;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12719; end if;
when s12720 => state := s12721; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12721 => 			--6
	if (mulfprdy = '1') then state := s12722;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12721; end if;
when s12722 => state := s12723; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12723 => 			--8
	if (mulfprdy = '1') then state := s12724;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12723; end if;
when s12724 => state := s12725; 	--9
	mulfpsclr <= '0';
when s12725 => state := s12726; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12726 => 			--11
	if (mulfprdy = '1') then state := s12727;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12726; end if;
when s12727 => state := s12728; 	--12
	mulfpsclr <= '0';
when s12728 => state := s12729; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12729 => 			--14
	if (addfprdy = '1') then state := s12730;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12729; end if;
when s12730 => state := s12731; 	--15
	addfpsclr <= '0';
when s12731 => state := s12732; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12732 => 			--17
	if (addfprdy = '1') then state := s12733;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12732; end if;
when s12733 => state := s12734; 	--18
	addfpsclr <= '0';
when s12734 => state := s12735; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12735 => 			--20
	if (addfprdy = '1') then state := s12736;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12735; end if;
when s12736 => state := s12737; 	--21
	addfpsclr <= '0';
when s12737 => state := s12738; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (634, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12738 => state := s12739; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1206, 12)); -- offset LSB 1158
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s12739 => state := s12740;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1207, 12)); -- offset MSB 1159
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12740 => state := s12741; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12741 => 			--4
	if (fixed2floatrdy = '1') then state := s12742;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12741; end if;
when s12742 => state := s12743; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12743 => 			--6
	if (mulfprdy = '1') then state := s12744;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12743; end if;
when s12744 => state := s12745; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12745 => 			--8
	if (mulfprdy = '1') then state := s12746;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12745; end if;
when s12746 => state := s12747; 	--9
	mulfpsclr <= '0';
when s12747 => state := s12748; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12748 => 			--11
	if (mulfprdy = '1') then state := s12749;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12748; end if;
when s12749 => state := s12750; 	--12
	mulfpsclr <= '0';
when s12750 => state := s12751; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12751 => 			--14
	if (addfprdy = '1') then state := s12752;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12751; end if;
when s12752 => state := s12753; 	--15
	addfpsclr <= '0';
when s12753 => state := s12754; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12754 => 			--17
	if (addfprdy = '1') then state := s12755;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12754; end if;
when s12755 => state := s12756; 	--18
	addfpsclr <= '0';
when s12756 => state := s12757; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12757 => 			--20
	if (addfprdy = '1') then state := s12758;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12757; end if;
when s12758 => state := s12759; 	--21
	addfpsclr <= '0';
when s12759 => state := s12760; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (635, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12760 => state := s12761; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1208, 12)); -- offset LSB 1160
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s12761 => state := s12762;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1209, 12)); -- offset MSB 1161
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12762 => state := s12763; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12763 => 			--4
	if (fixed2floatrdy = '1') then state := s12764;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12763; end if;
when s12764 => state := s12765; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12765 => 			--6
	if (mulfprdy = '1') then state := s12766;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12765; end if;
when s12766 => state := s12767; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12767 => 			--8
	if (mulfprdy = '1') then state := s12768;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12767; end if;
when s12768 => state := s12769; 	--9
	mulfpsclr <= '0';
when s12769 => state := s12770; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12770 => 			--11
	if (mulfprdy = '1') then state := s12771;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12770; end if;
when s12771 => state := s12772; 	--12
	mulfpsclr <= '0';
when s12772 => state := s12773; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12773 => 			--14
	if (addfprdy = '1') then state := s12774;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12773; end if;
when s12774 => state := s12775; 	--15
	addfpsclr <= '0';
when s12775 => state := s12776; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12776 => 			--17
	if (addfprdy = '1') then state := s12777;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12776; end if;
when s12777 => state := s12778; 	--18
	addfpsclr <= '0';
when s12778 => state := s12779; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12779 => 			--20
	if (addfprdy = '1') then state := s12780;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12779; end if;
when s12780 => state := s12781; 	--21
	addfpsclr <= '0';
when s12781 => state := s12782; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (636, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12782 => state := s12783; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1210, 12)); -- offset LSB 1162
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s12783 => state := s12784;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1211, 12)); -- offset MSB 1163
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12784 => state := s12785; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12785 => 			--4
	if (fixed2floatrdy = '1') then state := s12786;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12785; end if;
when s12786 => state := s12787; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12787 => 			--6
	if (mulfprdy = '1') then state := s12788;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12787; end if;
when s12788 => state := s12789; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12789 => 			--8
	if (mulfprdy = '1') then state := s12790;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12789; end if;
when s12790 => state := s12791; 	--9
	mulfpsclr <= '0';
when s12791 => state := s12792; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12792 => 			--11
	if (mulfprdy = '1') then state := s12793;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12792; end if;
when s12793 => state := s12794; 	--12
	mulfpsclr <= '0';
when s12794 => state := s12795; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12795 => 			--14
	if (addfprdy = '1') then state := s12796;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12795; end if;
when s12796 => state := s12797; 	--15
	addfpsclr <= '0';
when s12797 => state := s12798; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12798 => 			--17
	if (addfprdy = '1') then state := s12799;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12798; end if;
when s12799 => state := s12800; 	--18
	addfpsclr <= '0';
when s12800 => state := s12801; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12801 => 			--20
	if (addfprdy = '1') then state := s12802;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12801; end if;
when s12802 => state := s12803; 	--21
	addfpsclr <= '0';
when s12803 => state := s12804; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (637, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12804 => state := s12805; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1212, 12)); -- offset LSB 1164
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s12805 => state := s12806;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1213, 12)); -- offset MSB 1165
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12806 => state := s12807; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12807 => 			--4
	if (fixed2floatrdy = '1') then state := s12808;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12807; end if;
when s12808 => state := s12809; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12809 => 			--6
	if (mulfprdy = '1') then state := s12810;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12809; end if;
when s12810 => state := s12811; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12811 => 			--8
	if (mulfprdy = '1') then state := s12812;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12811; end if;
when s12812 => state := s12813; 	--9
	mulfpsclr <= '0';
when s12813 => state := s12814; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12814 => 			--11
	if (mulfprdy = '1') then state := s12815;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12814; end if;
when s12815 => state := s12816; 	--12
	mulfpsclr <= '0';
when s12816 => state := s12817; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12817 => 			--14
	if (addfprdy = '1') then state := s12818;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12817; end if;
when s12818 => state := s12819; 	--15
	addfpsclr <= '0';
when s12819 => state := s12820; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12820 => 			--17
	if (addfprdy = '1') then state := s12821;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12820; end if;
when s12821 => state := s12822; 	--18
	addfpsclr <= '0';
when s12822 => state := s12823; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12823 => 			--20
	if (addfprdy = '1') then state := s12824;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12823; end if;
when s12824 => state := s12825; 	--21
	addfpsclr <= '0';
when s12825 => state := s12826; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (638, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12826 => state := s12827; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1214, 12)); -- offset LSB 1166
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s12827 => state := s12828;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1215, 12)); -- offset MSB 1167
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12828 => state := s12829; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12829 => 			--4
	if (fixed2floatrdy = '1') then state := s12830;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12829; end if;
when s12830 => state := s12831; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12831 => 			--6
	if (mulfprdy = '1') then state := s12832;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12831; end if;
when s12832 => state := s12833; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12833 => 			--8
	if (mulfprdy = '1') then state := s12834;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12833; end if;
when s12834 => state := s12835; 	--9
	mulfpsclr <= '0';
when s12835 => state := s12836; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12836 => 			--11
	if (mulfprdy = '1') then state := s12837;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12836; end if;
when s12837 => state := s12838; 	--12
	mulfpsclr <= '0';
when s12838 => state := s12839; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12839 => 			--14
	if (addfprdy = '1') then state := s12840;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12839; end if;
when s12840 => state := s12841; 	--15
	addfpsclr <= '0';
when s12841 => state := s12842; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12842 => 			--17
	if (addfprdy = '1') then state := s12843;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12842; end if;
when s12843 => state := s12844; 	--18
	addfpsclr <= '0';
when s12844 => state := s12845; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12845 => 			--20
	if (addfprdy = '1') then state := s12846;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12845; end if;
when s12846 => state := s12847; 	--21
	addfpsclr <= '0';
when s12847 => state := s12848; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (639, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12848 => state := s12849; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1216, 12)); -- offset LSB 1168
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s12849 => state := s12850;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1217, 12)); -- offset MSB 1169
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12850 => state := s12851; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12851 => 			--4
	if (fixed2floatrdy = '1') then state := s12852;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12851; end if;
when s12852 => state := s12853; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12853 => 			--6
	if (mulfprdy = '1') then state := s12854;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12853; end if;
when s12854 => state := s12855; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12855 => 			--8
	if (mulfprdy = '1') then state := s12856;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12855; end if;
when s12856 => state := s12857; 	--9
	mulfpsclr <= '0';
when s12857 => state := s12858; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12858 => 			--11
	if (mulfprdy = '1') then state := s12859;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12858; end if;
when s12859 => state := s12860; 	--12
	mulfpsclr <= '0';
when s12860 => state := s12861; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12861 => 			--14
	if (addfprdy = '1') then state := s12862;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12861; end if;
when s12862 => state := s12863; 	--15
	addfpsclr <= '0';
when s12863 => state := s12864; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12864 => 			--17
	if (addfprdy = '1') then state := s12865;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12864; end if;
when s12865 => state := s12866; 	--18
	addfpsclr <= '0';
when s12866 => state := s12867; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12867 => 			--20
	if (addfprdy = '1') then state := s12868;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12867; end if;
when s12868 => state := s12869; 	--21
	addfpsclr <= '0';
when s12869 => state := s12870; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (640, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12870 => state := s12871; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1218, 12)); -- offset LSB 1170
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s12871 => state := s12872;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1219, 12)); -- offset MSB 1171
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12872 => state := s12873; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12873 => 			--4
	if (fixed2floatrdy = '1') then state := s12874;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12873; end if;
when s12874 => state := s12875; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12875 => 			--6
	if (mulfprdy = '1') then state := s12876;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12875; end if;
when s12876 => state := s12877; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12877 => 			--8
	if (mulfprdy = '1') then state := s12878;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12877; end if;
when s12878 => state := s12879; 	--9
	mulfpsclr <= '0';
when s12879 => state := s12880; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12880 => 			--11
	if (mulfprdy = '1') then state := s12881;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12880; end if;
when s12881 => state := s12882; 	--12
	mulfpsclr <= '0';
when s12882 => state := s12883; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12883 => 			--14
	if (addfprdy = '1') then state := s12884;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12883; end if;
when s12884 => state := s12885; 	--15
	addfpsclr <= '0';
when s12885 => state := s12886; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12886 => 			--17
	if (addfprdy = '1') then state := s12887;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12886; end if;
when s12887 => state := s12888; 	--18
	addfpsclr <= '0';
when s12888 => state := s12889; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12889 => 			--20
	if (addfprdy = '1') then state := s12890;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12889; end if;
when s12890 => state := s12891; 	--21
	addfpsclr <= '0';
when s12891 => state := s12892; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (641, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12892 => state := s12893; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1220, 12)); -- offset LSB 1172
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s12893 => state := s12894;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1221, 12)); -- offset MSB 1173
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12894 => state := s12895; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12895 => 			--4
	if (fixed2floatrdy = '1') then state := s12896;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12895; end if;
when s12896 => state := s12897; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12897 => 			--6
	if (mulfprdy = '1') then state := s12898;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12897; end if;
when s12898 => state := s12899; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12899 => 			--8
	if (mulfprdy = '1') then state := s12900;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12899; end if;
when s12900 => state := s12901; 	--9
	mulfpsclr <= '0';
when s12901 => state := s12902; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12902 => 			--11
	if (mulfprdy = '1') then state := s12903;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12902; end if;
when s12903 => state := s12904; 	--12
	mulfpsclr <= '0';
when s12904 => state := s12905; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12905 => 			--14
	if (addfprdy = '1') then state := s12906;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12905; end if;
when s12906 => state := s12907; 	--15
	addfpsclr <= '0';
when s12907 => state := s12908; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12908 => 			--17
	if (addfprdy = '1') then state := s12909;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12908; end if;
when s12909 => state := s12910; 	--18
	addfpsclr <= '0';
when s12910 => state := s12911; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12911 => 			--20
	if (addfprdy = '1') then state := s12912;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12911; end if;
when s12912 => state := s12913; 	--21
	addfpsclr <= '0';
when s12913 => state := s12914; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (642, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12914 => state := s12915; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1222, 12)); -- offset LSB 1174
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s12915 => state := s12916;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1223, 12)); -- offset MSB 1175
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12916 => state := s12917; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12917 => 			--4
	if (fixed2floatrdy = '1') then state := s12918;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12917; end if;
when s12918 => state := s12919; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12919 => 			--6
	if (mulfprdy = '1') then state := s12920;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12919; end if;
when s12920 => state := s12921; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12921 => 			--8
	if (mulfprdy = '1') then state := s12922;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12921; end if;
when s12922 => state := s12923; 	--9
	mulfpsclr <= '0';
when s12923 => state := s12924; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12924 => 			--11
	if (mulfprdy = '1') then state := s12925;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12924; end if;
when s12925 => state := s12926; 	--12
	mulfpsclr <= '0';
when s12926 => state := s12927; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12927 => 			--14
	if (addfprdy = '1') then state := s12928;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12927; end if;
when s12928 => state := s12929; 	--15
	addfpsclr <= '0';
when s12929 => state := s12930; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12930 => 			--17
	if (addfprdy = '1') then state := s12931;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12930; end if;
when s12931 => state := s12932; 	--18
	addfpsclr <= '0';
when s12932 => state := s12933; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12933 => 			--20
	if (addfprdy = '1') then state := s12934;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12933; end if;
when s12934 => state := s12935; 	--21
	addfpsclr <= '0';
when s12935 => state := s12936; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (643, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12936 => state := s12937; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1224, 12)); -- offset LSB 1176
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s12937 => state := s12938;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1225, 12)); -- offset MSB 1177
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12938 => state := s12939; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12939 => 			--4
	if (fixed2floatrdy = '1') then state := s12940;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12939; end if;
when s12940 => state := s12941; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12941 => 			--6
	if (mulfprdy = '1') then state := s12942;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12941; end if;
when s12942 => state := s12943; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12943 => 			--8
	if (mulfprdy = '1') then state := s12944;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12943; end if;
when s12944 => state := s12945; 	--9
	mulfpsclr <= '0';
when s12945 => state := s12946; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12946 => 			--11
	if (mulfprdy = '1') then state := s12947;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12946; end if;
when s12947 => state := s12948; 	--12
	mulfpsclr <= '0';
when s12948 => state := s12949; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12949 => 			--14
	if (addfprdy = '1') then state := s12950;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12949; end if;
when s12950 => state := s12951; 	--15
	addfpsclr <= '0';
when s12951 => state := s12952; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12952 => 			--17
	if (addfprdy = '1') then state := s12953;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12952; end if;
when s12953 => state := s12954; 	--18
	addfpsclr <= '0';
when s12954 => state := s12955; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12955 => 			--20
	if (addfprdy = '1') then state := s12956;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12955; end if;
when s12956 => state := s12957; 	--21
	addfpsclr <= '0';
when s12957 => state := s12958; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (644, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12958 => state := s12959; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1226, 12)); -- offset LSB 1178
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s12959 => state := s12960;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1227, 12)); -- offset MSB 1179
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12960 => state := s12961; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12961 => 			--4
	if (fixed2floatrdy = '1') then state := s12962;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12961; end if;
when s12962 => state := s12963; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12963 => 			--6
	if (mulfprdy = '1') then state := s12964;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12963; end if;
when s12964 => state := s12965; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12965 => 			--8
	if (mulfprdy = '1') then state := s12966;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12965; end if;
when s12966 => state := s12967; 	--9
	mulfpsclr <= '0';
when s12967 => state := s12968; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12968 => 			--11
	if (mulfprdy = '1') then state := s12969;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12968; end if;
when s12969 => state := s12970; 	--12
	mulfpsclr <= '0';
when s12970 => state := s12971; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12971 => 			--14
	if (addfprdy = '1') then state := s12972;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12971; end if;
when s12972 => state := s12973; 	--15
	addfpsclr <= '0';
when s12973 => state := s12974; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12974 => 			--17
	if (addfprdy = '1') then state := s12975;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12974; end if;
when s12975 => state := s12976; 	--18
	addfpsclr <= '0';
when s12976 => state := s12977; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12977 => 			--20
	if (addfprdy = '1') then state := s12978;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12977; end if;
when s12978 => state := s12979; 	--21
	addfpsclr <= '0';
when s12979 => state := s12980; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (645, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s12980 => state := s12981; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1228, 12)); -- offset LSB 1180
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s12981 => state := s12982;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1229, 12)); -- offset MSB 1181
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s12982 => state := s12983; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s12983 => 			--4
	if (fixed2floatrdy = '1') then state := s12984;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s12983; end if;
when s12984 => state := s12985; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s12985 => 			--6
	if (mulfprdy = '1') then state := s12986;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12985; end if;
when s12986 => state := s12987; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s12987 => 			--8
	if (mulfprdy = '1') then state := s12988;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12987; end if;
when s12988 => state := s12989; 	--9
	mulfpsclr <= '0';
when s12989 => state := s12990; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s12990 => 			--11
	if (mulfprdy = '1') then state := s12991;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s12990; end if;
when s12991 => state := s12992; 	--12
	mulfpsclr <= '0';
when s12992 => state := s12993; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s12993 => 			--14
	if (addfprdy = '1') then state := s12994;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12993; end if;
when s12994 => state := s12995; 	--15
	addfpsclr <= '0';
when s12995 => state := s12996; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s12996 => 			--17
	if (addfprdy = '1') then state := s12997;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12996; end if;
when s12997 => state := s12998; 	--18
	addfpsclr <= '0';
when s12998 => state := s12999; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s12999 => 			--20
	if (addfprdy = '1') then state := s13000;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s12999; end if;
when s13000 => state := s13001; 	--21
	addfpsclr <= '0';
when s13001 => state := s13002; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (646, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13002 => state := s13003; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1230, 12)); -- offset LSB 1182
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s13003 => state := s13004;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1231, 12)); -- offset MSB 1183
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13004 => state := s13005; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13005 => 			--4
	if (fixed2floatrdy = '1') then state := s13006;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13005; end if;
when s13006 => state := s13007; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13007 => 			--6
	if (mulfprdy = '1') then state := s13008;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13007; end if;
when s13008 => state := s13009; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13009 => 			--8
	if (mulfprdy = '1') then state := s13010;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13009; end if;
when s13010 => state := s13011; 	--9
	mulfpsclr <= '0';
when s13011 => state := s13012; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13012 => 			--11
	if (mulfprdy = '1') then state := s13013;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13012; end if;
when s13013 => state := s13014; 	--12
	mulfpsclr <= '0';
when s13014 => state := s13015; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13015 => 			--14
	if (addfprdy = '1') then state := s13016;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13015; end if;
when s13016 => state := s13017; 	--15
	addfpsclr <= '0';
when s13017 => state := s13018; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13018 => 			--17
	if (addfprdy = '1') then state := s13019;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13018; end if;
when s13019 => state := s13020; 	--18
	addfpsclr <= '0';
when s13020 => state := s13021; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13021 => 			--20
	if (addfprdy = '1') then state := s13022;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13021; end if;
when s13022 => state := s13023; 	--21
	addfpsclr <= '0';
when s13023 => state := s13024; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (647, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13024 => state := s13025; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1232, 12)); -- offset LSB 1184
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s13025 => state := s13026;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1233, 12)); -- offset MSB 1185
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13026 => state := s13027; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13027 => 			--4
	if (fixed2floatrdy = '1') then state := s13028;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13027; end if;
when s13028 => state := s13029; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13029 => 			--6
	if (mulfprdy = '1') then state := s13030;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13029; end if;
when s13030 => state := s13031; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13031 => 			--8
	if (mulfprdy = '1') then state := s13032;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13031; end if;
when s13032 => state := s13033; 	--9
	mulfpsclr <= '0';
when s13033 => state := s13034; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13034 => 			--11
	if (mulfprdy = '1') then state := s13035;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13034; end if;
when s13035 => state := s13036; 	--12
	mulfpsclr <= '0';
when s13036 => state := s13037; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13037 => 			--14
	if (addfprdy = '1') then state := s13038;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13037; end if;
when s13038 => state := s13039; 	--15
	addfpsclr <= '0';
when s13039 => state := s13040; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13040 => 			--17
	if (addfprdy = '1') then state := s13041;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13040; end if;
when s13041 => state := s13042; 	--18
	addfpsclr <= '0';
when s13042 => state := s13043; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13043 => 			--20
	if (addfprdy = '1') then state := s13044;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13043; end if;
when s13044 => state := s13045; 	--21
	addfpsclr <= '0';
when s13045 => state := s13046; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (648, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13046 => state := s13047; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1234, 12)); -- offset LSB 1186
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s13047 => state := s13048;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1235, 12)); -- offset MSB 1187
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13048 => state := s13049; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13049 => 			--4
	if (fixed2floatrdy = '1') then state := s13050;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13049; end if;
when s13050 => state := s13051; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13051 => 			--6
	if (mulfprdy = '1') then state := s13052;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13051; end if;
when s13052 => state := s13053; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13053 => 			--8
	if (mulfprdy = '1') then state := s13054;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13053; end if;
when s13054 => state := s13055; 	--9
	mulfpsclr <= '0';
when s13055 => state := s13056; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13056 => 			--11
	if (mulfprdy = '1') then state := s13057;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13056; end if;
when s13057 => state := s13058; 	--12
	mulfpsclr <= '0';
when s13058 => state := s13059; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13059 => 			--14
	if (addfprdy = '1') then state := s13060;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13059; end if;
when s13060 => state := s13061; 	--15
	addfpsclr <= '0';
when s13061 => state := s13062; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13062 => 			--17
	if (addfprdy = '1') then state := s13063;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13062; end if;
when s13063 => state := s13064; 	--18
	addfpsclr <= '0';
when s13064 => state := s13065; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13065 => 			--20
	if (addfprdy = '1') then state := s13066;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13065; end if;
when s13066 => state := s13067; 	--21
	addfpsclr <= '0';
when s13067 => state := s13068; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (649, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13068 => state := s13069; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1236, 12)); -- offset LSB 1188
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s13069 => state := s13070;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1237, 12)); -- offset MSB 1189
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13070 => state := s13071; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13071 => 			--4
	if (fixed2floatrdy = '1') then state := s13072;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13071; end if;
when s13072 => state := s13073; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13073 => 			--6
	if (mulfprdy = '1') then state := s13074;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13073; end if;
when s13074 => state := s13075; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13075 => 			--8
	if (mulfprdy = '1') then state := s13076;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13075; end if;
when s13076 => state := s13077; 	--9
	mulfpsclr <= '0';
when s13077 => state := s13078; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13078 => 			--11
	if (mulfprdy = '1') then state := s13079;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13078; end if;
when s13079 => state := s13080; 	--12
	mulfpsclr <= '0';
when s13080 => state := s13081; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13081 => 			--14
	if (addfprdy = '1') then state := s13082;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13081; end if;
when s13082 => state := s13083; 	--15
	addfpsclr <= '0';
when s13083 => state := s13084; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13084 => 			--17
	if (addfprdy = '1') then state := s13085;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13084; end if;
when s13085 => state := s13086; 	--18
	addfpsclr <= '0';
when s13086 => state := s13087; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13087 => 			--20
	if (addfprdy = '1') then state := s13088;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13087; end if;
when s13088 => state := s13089; 	--21
	addfpsclr <= '0';
when s13089 => state := s13090; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (650, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13090 => state := s13091; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1238, 12)); -- offset LSB 1190
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s13091 => state := s13092;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1239, 12)); -- offset MSB 1191
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13092 => state := s13093; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13093 => 			--4
	if (fixed2floatrdy = '1') then state := s13094;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13093; end if;
when s13094 => state := s13095; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13095 => 			--6
	if (mulfprdy = '1') then state := s13096;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13095; end if;
when s13096 => state := s13097; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13097 => 			--8
	if (mulfprdy = '1') then state := s13098;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13097; end if;
when s13098 => state := s13099; 	--9
	mulfpsclr <= '0';
when s13099 => state := s13100; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13100 => 			--11
	if (mulfprdy = '1') then state := s13101;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13100; end if;
when s13101 => state := s13102; 	--12
	mulfpsclr <= '0';
when s13102 => state := s13103; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13103 => 			--14
	if (addfprdy = '1') then state := s13104;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13103; end if;
when s13104 => state := s13105; 	--15
	addfpsclr <= '0';
when s13105 => state := s13106; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13106 => 			--17
	if (addfprdy = '1') then state := s13107;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13106; end if;
when s13107 => state := s13108; 	--18
	addfpsclr <= '0';
when s13108 => state := s13109; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13109 => 			--20
	if (addfprdy = '1') then state := s13110;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13109; end if;
when s13110 => state := s13111; 	--21
	addfpsclr <= '0';
when s13111 => state := s13112; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (651, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13112 => state := s13113; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1240, 12)); -- offset LSB 1192
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s13113 => state := s13114;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1241, 12)); -- offset MSB 1193
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13114 => state := s13115; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13115 => 			--4
	if (fixed2floatrdy = '1') then state := s13116;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13115; end if;
when s13116 => state := s13117; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13117 => 			--6
	if (mulfprdy = '1') then state := s13118;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13117; end if;
when s13118 => state := s13119; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13119 => 			--8
	if (mulfprdy = '1') then state := s13120;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13119; end if;
when s13120 => state := s13121; 	--9
	mulfpsclr <= '0';
when s13121 => state := s13122; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13122 => 			--11
	if (mulfprdy = '1') then state := s13123;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13122; end if;
when s13123 => state := s13124; 	--12
	mulfpsclr <= '0';
when s13124 => state := s13125; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13125 => 			--14
	if (addfprdy = '1') then state := s13126;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13125; end if;
when s13126 => state := s13127; 	--15
	addfpsclr <= '0';
when s13127 => state := s13128; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13128 => 			--17
	if (addfprdy = '1') then state := s13129;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13128; end if;
when s13129 => state := s13130; 	--18
	addfpsclr <= '0';
when s13130 => state := s13131; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13131 => 			--20
	if (addfprdy = '1') then state := s13132;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13131; end if;
when s13132 => state := s13133; 	--21
	addfpsclr <= '0';
when s13133 => state := s13134; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (652, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13134 => state := s13135; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1242, 12)); -- offset LSB 1194
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s13135 => state := s13136;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1243, 12)); -- offset MSB 1195
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13136 => state := s13137; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13137 => 			--4
	if (fixed2floatrdy = '1') then state := s13138;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13137; end if;
when s13138 => state := s13139; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13139 => 			--6
	if (mulfprdy = '1') then state := s13140;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13139; end if;
when s13140 => state := s13141; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13141 => 			--8
	if (mulfprdy = '1') then state := s13142;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13141; end if;
when s13142 => state := s13143; 	--9
	mulfpsclr <= '0';
when s13143 => state := s13144; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13144 => 			--11
	if (mulfprdy = '1') then state := s13145;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13144; end if;
when s13145 => state := s13146; 	--12
	mulfpsclr <= '0';
when s13146 => state := s13147; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13147 => 			--14
	if (addfprdy = '1') then state := s13148;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13147; end if;
when s13148 => state := s13149; 	--15
	addfpsclr <= '0';
when s13149 => state := s13150; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13150 => 			--17
	if (addfprdy = '1') then state := s13151;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13150; end if;
when s13151 => state := s13152; 	--18
	addfpsclr <= '0';
when s13152 => state := s13153; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13153 => 			--20
	if (addfprdy = '1') then state := s13154;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13153; end if;
when s13154 => state := s13155; 	--21
	addfpsclr <= '0';
when s13155 => state := s13156; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (653, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13156 => state := s13157; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1244, 12)); -- offset LSB 1196
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s13157 => state := s13158;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1245, 12)); -- offset MSB 1197
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13158 => state := s13159; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13159 => 			--4
	if (fixed2floatrdy = '1') then state := s13160;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13159; end if;
when s13160 => state := s13161; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13161 => 			--6
	if (mulfprdy = '1') then state := s13162;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13161; end if;
when s13162 => state := s13163; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13163 => 			--8
	if (mulfprdy = '1') then state := s13164;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13163; end if;
when s13164 => state := s13165; 	--9
	mulfpsclr <= '0';
when s13165 => state := s13166; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13166 => 			--11
	if (mulfprdy = '1') then state := s13167;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13166; end if;
when s13167 => state := s13168; 	--12
	mulfpsclr <= '0';
when s13168 => state := s13169; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13169 => 			--14
	if (addfprdy = '1') then state := s13170;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13169; end if;
when s13170 => state := s13171; 	--15
	addfpsclr <= '0';
when s13171 => state := s13172; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13172 => 			--17
	if (addfprdy = '1') then state := s13173;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13172; end if;
when s13173 => state := s13174; 	--18
	addfpsclr <= '0';
when s13174 => state := s13175; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13175 => 			--20
	if (addfprdy = '1') then state := s13176;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13175; end if;
when s13176 => state := s13177; 	--21
	addfpsclr <= '0';
when s13177 => state := s13178; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (654, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13178 => state := s13179; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1246, 12)); -- offset LSB 1198
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s13179 => state := s13180;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1247, 12)); -- offset MSB 1199
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13180 => state := s13181; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13181 => 			--4
	if (fixed2floatrdy = '1') then state := s13182;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13181; end if;
when s13182 => state := s13183; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13183 => 			--6
	if (mulfprdy = '1') then state := s13184;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13183; end if;
when s13184 => state := s13185; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13185 => 			--8
	if (mulfprdy = '1') then state := s13186;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13185; end if;
when s13186 => state := s13187; 	--9
	mulfpsclr <= '0';
when s13187 => state := s13188; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13188 => 			--11
	if (mulfprdy = '1') then state := s13189;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13188; end if;
when s13189 => state := s13190; 	--12
	mulfpsclr <= '0';
when s13190 => state := s13191; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13191 => 			--14
	if (addfprdy = '1') then state := s13192;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13191; end if;
when s13192 => state := s13193; 	--15
	addfpsclr <= '0';
when s13193 => state := s13194; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13194 => 			--17
	if (addfprdy = '1') then state := s13195;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13194; end if;
when s13195 => state := s13196; 	--18
	addfpsclr <= '0';
when s13196 => state := s13197; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13197 => 			--20
	if (addfprdy = '1') then state := s13198;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13197; end if;
when s13198 => state := s13199; 	--21
	addfpsclr <= '0';
when s13199 => state := s13200; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (655, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13200 => state := s13201; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1248, 12)); -- offset LSB 1200
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s13201 => state := s13202;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1249, 12)); -- offset MSB 1201
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13202 => state := s13203; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13203 => 			--4
	if (fixed2floatrdy = '1') then state := s13204;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13203; end if;
when s13204 => state := s13205; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13205 => 			--6
	if (mulfprdy = '1') then state := s13206;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13205; end if;
when s13206 => state := s13207; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13207 => 			--8
	if (mulfprdy = '1') then state := s13208;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13207; end if;
when s13208 => state := s13209; 	--9
	mulfpsclr <= '0';
when s13209 => state := s13210; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13210 => 			--11
	if (mulfprdy = '1') then state := s13211;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13210; end if;
when s13211 => state := s13212; 	--12
	mulfpsclr <= '0';
when s13212 => state := s13213; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13213 => 			--14
	if (addfprdy = '1') then state := s13214;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13213; end if;
when s13214 => state := s13215; 	--15
	addfpsclr <= '0';
when s13215 => state := s13216; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13216 => 			--17
	if (addfprdy = '1') then state := s13217;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13216; end if;
when s13217 => state := s13218; 	--18
	addfpsclr <= '0';
when s13218 => state := s13219; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13219 => 			--20
	if (addfprdy = '1') then state := s13220;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13219; end if;
when s13220 => state := s13221; 	--21
	addfpsclr <= '0';
when s13221 => state := s13222; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (656, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13222 => state := s13223; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1250, 12)); -- offset LSB 1202
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s13223 => state := s13224;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1251, 12)); -- offset MSB 1203
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13224 => state := s13225; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13225 => 			--4
	if (fixed2floatrdy = '1') then state := s13226;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13225; end if;
when s13226 => state := s13227; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13227 => 			--6
	if (mulfprdy = '1') then state := s13228;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13227; end if;
when s13228 => state := s13229; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13229 => 			--8
	if (mulfprdy = '1') then state := s13230;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13229; end if;
when s13230 => state := s13231; 	--9
	mulfpsclr <= '0';
when s13231 => state := s13232; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13232 => 			--11
	if (mulfprdy = '1') then state := s13233;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13232; end if;
when s13233 => state := s13234; 	--12
	mulfpsclr <= '0';
when s13234 => state := s13235; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13235 => 			--14
	if (addfprdy = '1') then state := s13236;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13235; end if;
when s13236 => state := s13237; 	--15
	addfpsclr <= '0';
when s13237 => state := s13238; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13238 => 			--17
	if (addfprdy = '1') then state := s13239;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13238; end if;
when s13239 => state := s13240; 	--18
	addfpsclr <= '0';
when s13240 => state := s13241; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13241 => 			--20
	if (addfprdy = '1') then state := s13242;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13241; end if;
when s13242 => state := s13243; 	--21
	addfpsclr <= '0';
when s13243 => state := s13244; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (657, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13244 => state := s13245; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1252, 12)); -- offset LSB 1204
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s13245 => state := s13246;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1253, 12)); -- offset MSB 1205
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13246 => state := s13247; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13247 => 			--4
	if (fixed2floatrdy = '1') then state := s13248;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13247; end if;
when s13248 => state := s13249; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13249 => 			--6
	if (mulfprdy = '1') then state := s13250;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13249; end if;
when s13250 => state := s13251; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13251 => 			--8
	if (mulfprdy = '1') then state := s13252;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13251; end if;
when s13252 => state := s13253; 	--9
	mulfpsclr <= '0';
when s13253 => state := s13254; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13254 => 			--11
	if (mulfprdy = '1') then state := s13255;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13254; end if;
when s13255 => state := s13256; 	--12
	mulfpsclr <= '0';
when s13256 => state := s13257; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13257 => 			--14
	if (addfprdy = '1') then state := s13258;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13257; end if;
when s13258 => state := s13259; 	--15
	addfpsclr <= '0';
when s13259 => state := s13260; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13260 => 			--17
	if (addfprdy = '1') then state := s13261;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13260; end if;
when s13261 => state := s13262; 	--18
	addfpsclr <= '0';
when s13262 => state := s13263; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13263 => 			--20
	if (addfprdy = '1') then state := s13264;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13263; end if;
when s13264 => state := s13265; 	--21
	addfpsclr <= '0';
when s13265 => state := s13266; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (658, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13266 => state := s13267; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1254, 12)); -- offset LSB 1206
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s13267 => state := s13268;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1255, 12)); -- offset MSB 1207
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13268 => state := s13269; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13269 => 			--4
	if (fixed2floatrdy = '1') then state := s13270;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13269; end if;
when s13270 => state := s13271; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13271 => 			--6
	if (mulfprdy = '1') then state := s13272;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13271; end if;
when s13272 => state := s13273; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13273 => 			--8
	if (mulfprdy = '1') then state := s13274;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13273; end if;
when s13274 => state := s13275; 	--9
	mulfpsclr <= '0';
when s13275 => state := s13276; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13276 => 			--11
	if (mulfprdy = '1') then state := s13277;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13276; end if;
when s13277 => state := s13278; 	--12
	mulfpsclr <= '0';
when s13278 => state := s13279; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13279 => 			--14
	if (addfprdy = '1') then state := s13280;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13279; end if;
when s13280 => state := s13281; 	--15
	addfpsclr <= '0';
when s13281 => state := s13282; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13282 => 			--17
	if (addfprdy = '1') then state := s13283;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13282; end if;
when s13283 => state := s13284; 	--18
	addfpsclr <= '0';
when s13284 => state := s13285; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13285 => 			--20
	if (addfprdy = '1') then state := s13286;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13285; end if;
when s13286 => state := s13287; 	--21
	addfpsclr <= '0';
when s13287 => state := s13288; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (659, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13288 => state := s13289; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1256, 12)); -- offset LSB 1208
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s13289 => state := s13290;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1257, 12)); -- offset MSB 1209
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13290 => state := s13291; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13291 => 			--4
	if (fixed2floatrdy = '1') then state := s13292;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13291; end if;
when s13292 => state := s13293; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13293 => 			--6
	if (mulfprdy = '1') then state := s13294;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13293; end if;
when s13294 => state := s13295; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13295 => 			--8
	if (mulfprdy = '1') then state := s13296;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13295; end if;
when s13296 => state := s13297; 	--9
	mulfpsclr <= '0';
when s13297 => state := s13298; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13298 => 			--11
	if (mulfprdy = '1') then state := s13299;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13298; end if;
when s13299 => state := s13300; 	--12
	mulfpsclr <= '0';
when s13300 => state := s13301; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13301 => 			--14
	if (addfprdy = '1') then state := s13302;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13301; end if;
when s13302 => state := s13303; 	--15
	addfpsclr <= '0';
when s13303 => state := s13304; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13304 => 			--17
	if (addfprdy = '1') then state := s13305;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13304; end if;
when s13305 => state := s13306; 	--18
	addfpsclr <= '0';
when s13306 => state := s13307; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13307 => 			--20
	if (addfprdy = '1') then state := s13308;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13307; end if;
when s13308 => state := s13309; 	--21
	addfpsclr <= '0';
when s13309 => state := s13310; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (660, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13310 => state := s13311; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1258, 12)); -- offset LSB 1210
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s13311 => state := s13312;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1259, 12)); -- offset MSB 1211
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13312 => state := s13313; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13313 => 			--4
	if (fixed2floatrdy = '1') then state := s13314;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13313; end if;
when s13314 => state := s13315; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13315 => 			--6
	if (mulfprdy = '1') then state := s13316;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13315; end if;
when s13316 => state := s13317; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13317 => 			--8
	if (mulfprdy = '1') then state := s13318;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13317; end if;
when s13318 => state := s13319; 	--9
	mulfpsclr <= '0';
when s13319 => state := s13320; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13320 => 			--11
	if (mulfprdy = '1') then state := s13321;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13320; end if;
when s13321 => state := s13322; 	--12
	mulfpsclr <= '0';
when s13322 => state := s13323; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13323 => 			--14
	if (addfprdy = '1') then state := s13324;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13323; end if;
when s13324 => state := s13325; 	--15
	addfpsclr <= '0';
when s13325 => state := s13326; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13326 => 			--17
	if (addfprdy = '1') then state := s13327;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13326; end if;
when s13327 => state := s13328; 	--18
	addfpsclr <= '0';
when s13328 => state := s13329; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13329 => 			--20
	if (addfprdy = '1') then state := s13330;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13329; end if;
when s13330 => state := s13331; 	--21
	addfpsclr <= '0';
when s13331 => state := s13332; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (661, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13332 => state := s13333; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1260, 12)); -- offset LSB 1212
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s13333 => state := s13334;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1261, 12)); -- offset MSB 1213
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13334 => state := s13335; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13335 => 			--4
	if (fixed2floatrdy = '1') then state := s13336;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13335; end if;
when s13336 => state := s13337; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13337 => 			--6
	if (mulfprdy = '1') then state := s13338;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13337; end if;
when s13338 => state := s13339; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13339 => 			--8
	if (mulfprdy = '1') then state := s13340;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13339; end if;
when s13340 => state := s13341; 	--9
	mulfpsclr <= '0';
when s13341 => state := s13342; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13342 => 			--11
	if (mulfprdy = '1') then state := s13343;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13342; end if;
when s13343 => state := s13344; 	--12
	mulfpsclr <= '0';
when s13344 => state := s13345; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13345 => 			--14
	if (addfprdy = '1') then state := s13346;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13345; end if;
when s13346 => state := s13347; 	--15
	addfpsclr <= '0';
when s13347 => state := s13348; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13348 => 			--17
	if (addfprdy = '1') then state := s13349;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13348; end if;
when s13349 => state := s13350; 	--18
	addfpsclr <= '0';
when s13350 => state := s13351; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13351 => 			--20
	if (addfprdy = '1') then state := s13352;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13351; end if;
when s13352 => state := s13353; 	--21
	addfpsclr <= '0';
when s13353 => state := s13354; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (662, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13354 => state := s13355; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1262, 12)); -- offset LSB 1214
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s13355 => state := s13356;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1263, 12)); -- offset MSB 1215
	addra <= std_logic_vector (to_unsigned (18, 10)); -- OCCrowI 18
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13356 => state := s13357; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13357 => 			--4
	if (fixed2floatrdy = '1') then state := s13358;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13357; end if;
when s13358 => state := s13359; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13359 => 			--6
	if (mulfprdy = '1') then state := s13360;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13359; end if;
when s13360 => state := s13361; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13361 => 			--8
	if (mulfprdy = '1') then state := s13362;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13361; end if;
when s13362 => state := s13363; 	--9
	mulfpsclr <= '0';
when s13363 => state := s13364; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13364 => 			--11
	if (mulfprdy = '1') then state := s13365;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13364; end if;
when s13365 => state := s13366; 	--12
	mulfpsclr <= '0';
when s13366 => state := s13367; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13367 => 			--14
	if (addfprdy = '1') then state := s13368;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13367; end if;
when s13368 => state := s13369; 	--15
	addfpsclr <= '0';
when s13369 => state := s13370; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13370 => 			--17
	if (addfprdy = '1') then state := s13371;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13370; end if;
when s13371 => state := s13372; 	--18
	addfpsclr <= '0';
when s13372 => state := s13373; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13373 => 			--20
	if (addfprdy = '1') then state := s13374;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13373; end if;
when s13374 => state := s13375; 	--21
	addfpsclr <= '0';
when s13375 => state := s13376; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (663, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13376 => state := s13377; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1264, 12)); -- offset LSB 1216
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s13377 => state := s13378;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1265, 12)); -- offset MSB 1217
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13378 => state := s13379; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13379 => 			--4
	if (fixed2floatrdy = '1') then state := s13380;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13379; end if;
when s13380 => state := s13381; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13381 => 			--6
	if (mulfprdy = '1') then state := s13382;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13381; end if;
when s13382 => state := s13383; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13383 => 			--8
	if (mulfprdy = '1') then state := s13384;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13383; end if;
when s13384 => state := s13385; 	--9
	mulfpsclr <= '0';
when s13385 => state := s13386; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13386 => 			--11
	if (mulfprdy = '1') then state := s13387;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13386; end if;
when s13387 => state := s13388; 	--12
	mulfpsclr <= '0';
when s13388 => state := s13389; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13389 => 			--14
	if (addfprdy = '1') then state := s13390;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13389; end if;
when s13390 => state := s13391; 	--15
	addfpsclr <= '0';
when s13391 => state := s13392; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13392 => 			--17
	if (addfprdy = '1') then state := s13393;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13392; end if;
when s13393 => state := s13394; 	--18
	addfpsclr <= '0';
when s13394 => state := s13395; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13395 => 			--20
	if (addfprdy = '1') then state := s13396;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13395; end if;
when s13396 => state := s13397; 	--21
	addfpsclr <= '0';
when s13397 => state := s13398; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (664, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13398 => state := s13399; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1266, 12)); -- offset LSB 1218
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s13399 => state := s13400;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1267, 12)); -- offset MSB 1219
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13400 => state := s13401; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13401 => 			--4
	if (fixed2floatrdy = '1') then state := s13402;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13401; end if;
when s13402 => state := s13403; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13403 => 			--6
	if (mulfprdy = '1') then state := s13404;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13403; end if;
when s13404 => state := s13405; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13405 => 			--8
	if (mulfprdy = '1') then state := s13406;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13405; end if;
when s13406 => state := s13407; 	--9
	mulfpsclr <= '0';
when s13407 => state := s13408; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13408 => 			--11
	if (mulfprdy = '1') then state := s13409;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13408; end if;
when s13409 => state := s13410; 	--12
	mulfpsclr <= '0';
when s13410 => state := s13411; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13411 => 			--14
	if (addfprdy = '1') then state := s13412;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13411; end if;
when s13412 => state := s13413; 	--15
	addfpsclr <= '0';
when s13413 => state := s13414; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13414 => 			--17
	if (addfprdy = '1') then state := s13415;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13414; end if;
when s13415 => state := s13416; 	--18
	addfpsclr <= '0';
when s13416 => state := s13417; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13417 => 			--20
	if (addfprdy = '1') then state := s13418;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13417; end if;
when s13418 => state := s13419; 	--21
	addfpsclr <= '0';
when s13419 => state := s13420; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (665, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13420 => state := s13421; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1268, 12)); -- offset LSB 1220
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s13421 => state := s13422;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1269, 12)); -- offset MSB 1221
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13422 => state := s13423; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13423 => 			--4
	if (fixed2floatrdy = '1') then state := s13424;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13423; end if;
when s13424 => state := s13425; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13425 => 			--6
	if (mulfprdy = '1') then state := s13426;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13425; end if;
when s13426 => state := s13427; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13427 => 			--8
	if (mulfprdy = '1') then state := s13428;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13427; end if;
when s13428 => state := s13429; 	--9
	mulfpsclr <= '0';
when s13429 => state := s13430; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13430 => 			--11
	if (mulfprdy = '1') then state := s13431;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13430; end if;
when s13431 => state := s13432; 	--12
	mulfpsclr <= '0';
when s13432 => state := s13433; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13433 => 			--14
	if (addfprdy = '1') then state := s13434;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13433; end if;
when s13434 => state := s13435; 	--15
	addfpsclr <= '0';
when s13435 => state := s13436; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13436 => 			--17
	if (addfprdy = '1') then state := s13437;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13436; end if;
when s13437 => state := s13438; 	--18
	addfpsclr <= '0';
when s13438 => state := s13439; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13439 => 			--20
	if (addfprdy = '1') then state := s13440;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13439; end if;
when s13440 => state := s13441; 	--21
	addfpsclr <= '0';
when s13441 => state := s13442; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (666, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13442 => state := s13443; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1270, 12)); -- offset LSB 1222
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s13443 => state := s13444;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1271, 12)); -- offset MSB 1223
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13444 => state := s13445; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13445 => 			--4
	if (fixed2floatrdy = '1') then state := s13446;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13445; end if;
when s13446 => state := s13447; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13447 => 			--6
	if (mulfprdy = '1') then state := s13448;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13447; end if;
when s13448 => state := s13449; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13449 => 			--8
	if (mulfprdy = '1') then state := s13450;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13449; end if;
when s13450 => state := s13451; 	--9
	mulfpsclr <= '0';
when s13451 => state := s13452; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13452 => 			--11
	if (mulfprdy = '1') then state := s13453;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13452; end if;
when s13453 => state := s13454; 	--12
	mulfpsclr <= '0';
when s13454 => state := s13455; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13455 => 			--14
	if (addfprdy = '1') then state := s13456;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13455; end if;
when s13456 => state := s13457; 	--15
	addfpsclr <= '0';
when s13457 => state := s13458; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13458 => 			--17
	if (addfprdy = '1') then state := s13459;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13458; end if;
when s13459 => state := s13460; 	--18
	addfpsclr <= '0';
when s13460 => state := s13461; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13461 => 			--20
	if (addfprdy = '1') then state := s13462;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13461; end if;
when s13462 => state := s13463; 	--21
	addfpsclr <= '0';
when s13463 => state := s13464; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (667, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13464 => state := s13465; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1272, 12)); -- offset LSB 1224
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s13465 => state := s13466;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1273, 12)); -- offset MSB 1225
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13466 => state := s13467; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13467 => 			--4
	if (fixed2floatrdy = '1') then state := s13468;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13467; end if;
when s13468 => state := s13469; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13469 => 			--6
	if (mulfprdy = '1') then state := s13470;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13469; end if;
when s13470 => state := s13471; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13471 => 			--8
	if (mulfprdy = '1') then state := s13472;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13471; end if;
when s13472 => state := s13473; 	--9
	mulfpsclr <= '0';
when s13473 => state := s13474; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13474 => 			--11
	if (mulfprdy = '1') then state := s13475;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13474; end if;
when s13475 => state := s13476; 	--12
	mulfpsclr <= '0';
when s13476 => state := s13477; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13477 => 			--14
	if (addfprdy = '1') then state := s13478;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13477; end if;
when s13478 => state := s13479; 	--15
	addfpsclr <= '0';
when s13479 => state := s13480; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13480 => 			--17
	if (addfprdy = '1') then state := s13481;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13480; end if;
when s13481 => state := s13482; 	--18
	addfpsclr <= '0';
when s13482 => state := s13483; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13483 => 			--20
	if (addfprdy = '1') then state := s13484;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13483; end if;
when s13484 => state := s13485; 	--21
	addfpsclr <= '0';
when s13485 => state := s13486; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (668, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13486 => state := s13487; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1274, 12)); -- offset LSB 1226
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s13487 => state := s13488;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1275, 12)); -- offset MSB 1227
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13488 => state := s13489; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13489 => 			--4
	if (fixed2floatrdy = '1') then state := s13490;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13489; end if;
when s13490 => state := s13491; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13491 => 			--6
	if (mulfprdy = '1') then state := s13492;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13491; end if;
when s13492 => state := s13493; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13493 => 			--8
	if (mulfprdy = '1') then state := s13494;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13493; end if;
when s13494 => state := s13495; 	--9
	mulfpsclr <= '0';
when s13495 => state := s13496; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13496 => 			--11
	if (mulfprdy = '1') then state := s13497;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13496; end if;
when s13497 => state := s13498; 	--12
	mulfpsclr <= '0';
when s13498 => state := s13499; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13499 => 			--14
	if (addfprdy = '1') then state := s13500;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13499; end if;
when s13500 => state := s13501; 	--15
	addfpsclr <= '0';
when s13501 => state := s13502; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13502 => 			--17
	if (addfprdy = '1') then state := s13503;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13502; end if;
when s13503 => state := s13504; 	--18
	addfpsclr <= '0';
when s13504 => state := s13505; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13505 => 			--20
	if (addfprdy = '1') then state := s13506;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13505; end if;
when s13506 => state := s13507; 	--21
	addfpsclr <= '0';
when s13507 => state := s13508; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (669, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13508 => state := s13509; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1276, 12)); -- offset LSB 1228
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s13509 => state := s13510;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1277, 12)); -- offset MSB 1229
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13510 => state := s13511; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13511 => 			--4
	if (fixed2floatrdy = '1') then state := s13512;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13511; end if;
when s13512 => state := s13513; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13513 => 			--6
	if (mulfprdy = '1') then state := s13514;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13513; end if;
when s13514 => state := s13515; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13515 => 			--8
	if (mulfprdy = '1') then state := s13516;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13515; end if;
when s13516 => state := s13517; 	--9
	mulfpsclr <= '0';
when s13517 => state := s13518; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13518 => 			--11
	if (mulfprdy = '1') then state := s13519;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13518; end if;
when s13519 => state := s13520; 	--12
	mulfpsclr <= '0';
when s13520 => state := s13521; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13521 => 			--14
	if (addfprdy = '1') then state := s13522;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13521; end if;
when s13522 => state := s13523; 	--15
	addfpsclr <= '0';
when s13523 => state := s13524; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13524 => 			--17
	if (addfprdy = '1') then state := s13525;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13524; end if;
when s13525 => state := s13526; 	--18
	addfpsclr <= '0';
when s13526 => state := s13527; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13527 => 			--20
	if (addfprdy = '1') then state := s13528;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13527; end if;
when s13528 => state := s13529; 	--21
	addfpsclr <= '0';
when s13529 => state := s13530; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (670, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13530 => state := s13531; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1278, 12)); -- offset LSB 1230
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s13531 => state := s13532;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1279, 12)); -- offset MSB 1231
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13532 => state := s13533; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13533 => 			--4
	if (fixed2floatrdy = '1') then state := s13534;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13533; end if;
when s13534 => state := s13535; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13535 => 			--6
	if (mulfprdy = '1') then state := s13536;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13535; end if;
when s13536 => state := s13537; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13537 => 			--8
	if (mulfprdy = '1') then state := s13538;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13537; end if;
when s13538 => state := s13539; 	--9
	mulfpsclr <= '0';
when s13539 => state := s13540; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13540 => 			--11
	if (mulfprdy = '1') then state := s13541;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13540; end if;
when s13541 => state := s13542; 	--12
	mulfpsclr <= '0';
when s13542 => state := s13543; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13543 => 			--14
	if (addfprdy = '1') then state := s13544;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13543; end if;
when s13544 => state := s13545; 	--15
	addfpsclr <= '0';
when s13545 => state := s13546; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13546 => 			--17
	if (addfprdy = '1') then state := s13547;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13546; end if;
when s13547 => state := s13548; 	--18
	addfpsclr <= '0';
when s13548 => state := s13549; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13549 => 			--20
	if (addfprdy = '1') then state := s13550;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13549; end if;
when s13550 => state := s13551; 	--21
	addfpsclr <= '0';
when s13551 => state := s13552; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (671, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13552 => state := s13553; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1280, 12)); -- offset LSB 1232
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s13553 => state := s13554;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1281, 12)); -- offset MSB 1233
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13554 => state := s13555; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13555 => 			--4
	if (fixed2floatrdy = '1') then state := s13556;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13555; end if;
when s13556 => state := s13557; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13557 => 			--6
	if (mulfprdy = '1') then state := s13558;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13557; end if;
when s13558 => state := s13559; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13559 => 			--8
	if (mulfprdy = '1') then state := s13560;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13559; end if;
when s13560 => state := s13561; 	--9
	mulfpsclr <= '0';
when s13561 => state := s13562; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13562 => 			--11
	if (mulfprdy = '1') then state := s13563;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13562; end if;
when s13563 => state := s13564; 	--12
	mulfpsclr <= '0';
when s13564 => state := s13565; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13565 => 			--14
	if (addfprdy = '1') then state := s13566;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13565; end if;
when s13566 => state := s13567; 	--15
	addfpsclr <= '0';
when s13567 => state := s13568; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13568 => 			--17
	if (addfprdy = '1') then state := s13569;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13568; end if;
when s13569 => state := s13570; 	--18
	addfpsclr <= '0';
when s13570 => state := s13571; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13571 => 			--20
	if (addfprdy = '1') then state := s13572;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13571; end if;
when s13572 => state := s13573; 	--21
	addfpsclr <= '0';
when s13573 => state := s13574; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (672, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13574 => state := s13575; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1282, 12)); -- offset LSB 1234
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s13575 => state := s13576;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1283, 12)); -- offset MSB 1235
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13576 => state := s13577; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13577 => 			--4
	if (fixed2floatrdy = '1') then state := s13578;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13577; end if;
when s13578 => state := s13579; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13579 => 			--6
	if (mulfprdy = '1') then state := s13580;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13579; end if;
when s13580 => state := s13581; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13581 => 			--8
	if (mulfprdy = '1') then state := s13582;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13581; end if;
when s13582 => state := s13583; 	--9
	mulfpsclr <= '0';
when s13583 => state := s13584; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13584 => 			--11
	if (mulfprdy = '1') then state := s13585;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13584; end if;
when s13585 => state := s13586; 	--12
	mulfpsclr <= '0';
when s13586 => state := s13587; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13587 => 			--14
	if (addfprdy = '1') then state := s13588;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13587; end if;
when s13588 => state := s13589; 	--15
	addfpsclr <= '0';
when s13589 => state := s13590; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13590 => 			--17
	if (addfprdy = '1') then state := s13591;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13590; end if;
when s13591 => state := s13592; 	--18
	addfpsclr <= '0';
when s13592 => state := s13593; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13593 => 			--20
	if (addfprdy = '1') then state := s13594;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13593; end if;
when s13594 => state := s13595; 	--21
	addfpsclr <= '0';
when s13595 => state := s13596; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (673, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13596 => state := s13597; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1284, 12)); -- offset LSB 1236
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s13597 => state := s13598;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1285, 12)); -- offset MSB 1237
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13598 => state := s13599; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13599 => 			--4
	if (fixed2floatrdy = '1') then state := s13600;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13599; end if;
when s13600 => state := s13601; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13601 => 			--6
	if (mulfprdy = '1') then state := s13602;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13601; end if;
when s13602 => state := s13603; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13603 => 			--8
	if (mulfprdy = '1') then state := s13604;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13603; end if;
when s13604 => state := s13605; 	--9
	mulfpsclr <= '0';
when s13605 => state := s13606; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13606 => 			--11
	if (mulfprdy = '1') then state := s13607;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13606; end if;
when s13607 => state := s13608; 	--12
	mulfpsclr <= '0';
when s13608 => state := s13609; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13609 => 			--14
	if (addfprdy = '1') then state := s13610;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13609; end if;
when s13610 => state := s13611; 	--15
	addfpsclr <= '0';
when s13611 => state := s13612; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13612 => 			--17
	if (addfprdy = '1') then state := s13613;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13612; end if;
when s13613 => state := s13614; 	--18
	addfpsclr <= '0';
when s13614 => state := s13615; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13615 => 			--20
	if (addfprdy = '1') then state := s13616;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13615; end if;
when s13616 => state := s13617; 	--21
	addfpsclr <= '0';
when s13617 => state := s13618; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (674, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13618 => state := s13619; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1286, 12)); -- offset LSB 1238
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s13619 => state := s13620;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1287, 12)); -- offset MSB 1239
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13620 => state := s13621; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13621 => 			--4
	if (fixed2floatrdy = '1') then state := s13622;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13621; end if;
when s13622 => state := s13623; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13623 => 			--6
	if (mulfprdy = '1') then state := s13624;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13623; end if;
when s13624 => state := s13625; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13625 => 			--8
	if (mulfprdy = '1') then state := s13626;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13625; end if;
when s13626 => state := s13627; 	--9
	mulfpsclr <= '0';
when s13627 => state := s13628; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13628 => 			--11
	if (mulfprdy = '1') then state := s13629;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13628; end if;
when s13629 => state := s13630; 	--12
	mulfpsclr <= '0';
when s13630 => state := s13631; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13631 => 			--14
	if (addfprdy = '1') then state := s13632;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13631; end if;
when s13632 => state := s13633; 	--15
	addfpsclr <= '0';
when s13633 => state := s13634; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13634 => 			--17
	if (addfprdy = '1') then state := s13635;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13634; end if;
when s13635 => state := s13636; 	--18
	addfpsclr <= '0';
when s13636 => state := s13637; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13637 => 			--20
	if (addfprdy = '1') then state := s13638;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13637; end if;
when s13638 => state := s13639; 	--21
	addfpsclr <= '0';
when s13639 => state := s13640; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (675, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13640 => state := s13641; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1288, 12)); -- offset LSB 1240
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s13641 => state := s13642;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1289, 12)); -- offset MSB 1241
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13642 => state := s13643; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13643 => 			--4
	if (fixed2floatrdy = '1') then state := s13644;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13643; end if;
when s13644 => state := s13645; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13645 => 			--6
	if (mulfprdy = '1') then state := s13646;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13645; end if;
when s13646 => state := s13647; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13647 => 			--8
	if (mulfprdy = '1') then state := s13648;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13647; end if;
when s13648 => state := s13649; 	--9
	mulfpsclr <= '0';
when s13649 => state := s13650; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13650 => 			--11
	if (mulfprdy = '1') then state := s13651;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13650; end if;
when s13651 => state := s13652; 	--12
	mulfpsclr <= '0';
when s13652 => state := s13653; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13653 => 			--14
	if (addfprdy = '1') then state := s13654;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13653; end if;
when s13654 => state := s13655; 	--15
	addfpsclr <= '0';
when s13655 => state := s13656; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13656 => 			--17
	if (addfprdy = '1') then state := s13657;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13656; end if;
when s13657 => state := s13658; 	--18
	addfpsclr <= '0';
when s13658 => state := s13659; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13659 => 			--20
	if (addfprdy = '1') then state := s13660;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13659; end if;
when s13660 => state := s13661; 	--21
	addfpsclr <= '0';
when s13661 => state := s13662; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (676, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13662 => state := s13663; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1290, 12)); -- offset LSB 1242
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s13663 => state := s13664;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1291, 12)); -- offset MSB 1243
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13664 => state := s13665; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13665 => 			--4
	if (fixed2floatrdy = '1') then state := s13666;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13665; end if;
when s13666 => state := s13667; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13667 => 			--6
	if (mulfprdy = '1') then state := s13668;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13667; end if;
when s13668 => state := s13669; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13669 => 			--8
	if (mulfprdy = '1') then state := s13670;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13669; end if;
when s13670 => state := s13671; 	--9
	mulfpsclr <= '0';
when s13671 => state := s13672; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13672 => 			--11
	if (mulfprdy = '1') then state := s13673;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13672; end if;
when s13673 => state := s13674; 	--12
	mulfpsclr <= '0';
when s13674 => state := s13675; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13675 => 			--14
	if (addfprdy = '1') then state := s13676;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13675; end if;
when s13676 => state := s13677; 	--15
	addfpsclr <= '0';
when s13677 => state := s13678; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13678 => 			--17
	if (addfprdy = '1') then state := s13679;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13678; end if;
when s13679 => state := s13680; 	--18
	addfpsclr <= '0';
when s13680 => state := s13681; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13681 => 			--20
	if (addfprdy = '1') then state := s13682;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13681; end if;
when s13682 => state := s13683; 	--21
	addfpsclr <= '0';
when s13683 => state := s13684; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (677, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13684 => state := s13685; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1292, 12)); -- offset LSB 1244
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s13685 => state := s13686;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1293, 12)); -- offset MSB 1245
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13686 => state := s13687; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13687 => 			--4
	if (fixed2floatrdy = '1') then state := s13688;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13687; end if;
when s13688 => state := s13689; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13689 => 			--6
	if (mulfprdy = '1') then state := s13690;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13689; end if;
when s13690 => state := s13691; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13691 => 			--8
	if (mulfprdy = '1') then state := s13692;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13691; end if;
when s13692 => state := s13693; 	--9
	mulfpsclr <= '0';
when s13693 => state := s13694; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13694 => 			--11
	if (mulfprdy = '1') then state := s13695;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13694; end if;
when s13695 => state := s13696; 	--12
	mulfpsclr <= '0';
when s13696 => state := s13697; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13697 => 			--14
	if (addfprdy = '1') then state := s13698;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13697; end if;
when s13698 => state := s13699; 	--15
	addfpsclr <= '0';
when s13699 => state := s13700; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13700 => 			--17
	if (addfprdy = '1') then state := s13701;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13700; end if;
when s13701 => state := s13702; 	--18
	addfpsclr <= '0';
when s13702 => state := s13703; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13703 => 			--20
	if (addfprdy = '1') then state := s13704;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13703; end if;
when s13704 => state := s13705; 	--21
	addfpsclr <= '0';
when s13705 => state := s13706; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (678, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13706 => state := s13707; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1294, 12)); -- offset LSB 1246
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s13707 => state := s13708;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1295, 12)); -- offset MSB 1247
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13708 => state := s13709; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13709 => 			--4
	if (fixed2floatrdy = '1') then state := s13710;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13709; end if;
when s13710 => state := s13711; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13711 => 			--6
	if (mulfprdy = '1') then state := s13712;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13711; end if;
when s13712 => state := s13713; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13713 => 			--8
	if (mulfprdy = '1') then state := s13714;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13713; end if;
when s13714 => state := s13715; 	--9
	mulfpsclr <= '0';
when s13715 => state := s13716; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13716 => 			--11
	if (mulfprdy = '1') then state := s13717;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13716; end if;
when s13717 => state := s13718; 	--12
	mulfpsclr <= '0';
when s13718 => state := s13719; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13719 => 			--14
	if (addfprdy = '1') then state := s13720;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13719; end if;
when s13720 => state := s13721; 	--15
	addfpsclr <= '0';
when s13721 => state := s13722; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13722 => 			--17
	if (addfprdy = '1') then state := s13723;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13722; end if;
when s13723 => state := s13724; 	--18
	addfpsclr <= '0';
when s13724 => state := s13725; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13725 => 			--20
	if (addfprdy = '1') then state := s13726;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13725; end if;
when s13726 => state := s13727; 	--21
	addfpsclr <= '0';
when s13727 => state := s13728; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (679, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13728 => state := s13729; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1296, 12)); -- offset LSB 1248
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s13729 => state := s13730;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1297, 12)); -- offset MSB 1249
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13730 => state := s13731; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13731 => 			--4
	if (fixed2floatrdy = '1') then state := s13732;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13731; end if;
when s13732 => state := s13733; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13733 => 			--6
	if (mulfprdy = '1') then state := s13734;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13733; end if;
when s13734 => state := s13735; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13735 => 			--8
	if (mulfprdy = '1') then state := s13736;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13735; end if;
when s13736 => state := s13737; 	--9
	mulfpsclr <= '0';
when s13737 => state := s13738; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13738 => 			--11
	if (mulfprdy = '1') then state := s13739;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13738; end if;
when s13739 => state := s13740; 	--12
	mulfpsclr <= '0';
when s13740 => state := s13741; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13741 => 			--14
	if (addfprdy = '1') then state := s13742;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13741; end if;
when s13742 => state := s13743; 	--15
	addfpsclr <= '0';
when s13743 => state := s13744; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13744 => 			--17
	if (addfprdy = '1') then state := s13745;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13744; end if;
when s13745 => state := s13746; 	--18
	addfpsclr <= '0';
when s13746 => state := s13747; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13747 => 			--20
	if (addfprdy = '1') then state := s13748;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13747; end if;
when s13748 => state := s13749; 	--21
	addfpsclr <= '0';
when s13749 => state := s13750; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (680, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13750 => state := s13751; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1298, 12)); -- offset LSB 1250
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s13751 => state := s13752;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1299, 12)); -- offset MSB 1251
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13752 => state := s13753; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13753 => 			--4
	if (fixed2floatrdy = '1') then state := s13754;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13753; end if;
when s13754 => state := s13755; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13755 => 			--6
	if (mulfprdy = '1') then state := s13756;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13755; end if;
when s13756 => state := s13757; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13757 => 			--8
	if (mulfprdy = '1') then state := s13758;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13757; end if;
when s13758 => state := s13759; 	--9
	mulfpsclr <= '0';
when s13759 => state := s13760; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13760 => 			--11
	if (mulfprdy = '1') then state := s13761;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13760; end if;
when s13761 => state := s13762; 	--12
	mulfpsclr <= '0';
when s13762 => state := s13763; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13763 => 			--14
	if (addfprdy = '1') then state := s13764;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13763; end if;
when s13764 => state := s13765; 	--15
	addfpsclr <= '0';
when s13765 => state := s13766; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13766 => 			--17
	if (addfprdy = '1') then state := s13767;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13766; end if;
when s13767 => state := s13768; 	--18
	addfpsclr <= '0';
when s13768 => state := s13769; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13769 => 			--20
	if (addfprdy = '1') then state := s13770;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13769; end if;
when s13770 => state := s13771; 	--21
	addfpsclr <= '0';
when s13771 => state := s13772; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (681, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13772 => state := s13773; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1300, 12)); -- offset LSB 1252
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s13773 => state := s13774;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1301, 12)); -- offset MSB 1253
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13774 => state := s13775; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13775 => 			--4
	if (fixed2floatrdy = '1') then state := s13776;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13775; end if;
when s13776 => state := s13777; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13777 => 			--6
	if (mulfprdy = '1') then state := s13778;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13777; end if;
when s13778 => state := s13779; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13779 => 			--8
	if (mulfprdy = '1') then state := s13780;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13779; end if;
when s13780 => state := s13781; 	--9
	mulfpsclr <= '0';
when s13781 => state := s13782; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13782 => 			--11
	if (mulfprdy = '1') then state := s13783;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13782; end if;
when s13783 => state := s13784; 	--12
	mulfpsclr <= '0';
when s13784 => state := s13785; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13785 => 			--14
	if (addfprdy = '1') then state := s13786;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13785; end if;
when s13786 => state := s13787; 	--15
	addfpsclr <= '0';
when s13787 => state := s13788; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13788 => 			--17
	if (addfprdy = '1') then state := s13789;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13788; end if;
when s13789 => state := s13790; 	--18
	addfpsclr <= '0';
when s13790 => state := s13791; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13791 => 			--20
	if (addfprdy = '1') then state := s13792;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13791; end if;
when s13792 => state := s13793; 	--21
	addfpsclr <= '0';
when s13793 => state := s13794; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (682, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13794 => state := s13795; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1302, 12)); -- offset LSB 1254
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s13795 => state := s13796;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1303, 12)); -- offset MSB 1255
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13796 => state := s13797; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13797 => 			--4
	if (fixed2floatrdy = '1') then state := s13798;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13797; end if;
when s13798 => state := s13799; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13799 => 			--6
	if (mulfprdy = '1') then state := s13800;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13799; end if;
when s13800 => state := s13801; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13801 => 			--8
	if (mulfprdy = '1') then state := s13802;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13801; end if;
when s13802 => state := s13803; 	--9
	mulfpsclr <= '0';
when s13803 => state := s13804; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13804 => 			--11
	if (mulfprdy = '1') then state := s13805;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13804; end if;
when s13805 => state := s13806; 	--12
	mulfpsclr <= '0';
when s13806 => state := s13807; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13807 => 			--14
	if (addfprdy = '1') then state := s13808;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13807; end if;
when s13808 => state := s13809; 	--15
	addfpsclr <= '0';
when s13809 => state := s13810; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13810 => 			--17
	if (addfprdy = '1') then state := s13811;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13810; end if;
when s13811 => state := s13812; 	--18
	addfpsclr <= '0';
when s13812 => state := s13813; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13813 => 			--20
	if (addfprdy = '1') then state := s13814;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13813; end if;
when s13814 => state := s13815; 	--21
	addfpsclr <= '0';
when s13815 => state := s13816; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (683, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13816 => state := s13817; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1304, 12)); -- offset LSB 1256
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s13817 => state := s13818;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1305, 12)); -- offset MSB 1257
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13818 => state := s13819; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13819 => 			--4
	if (fixed2floatrdy = '1') then state := s13820;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13819; end if;
when s13820 => state := s13821; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13821 => 			--6
	if (mulfprdy = '1') then state := s13822;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13821; end if;
when s13822 => state := s13823; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13823 => 			--8
	if (mulfprdy = '1') then state := s13824;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13823; end if;
when s13824 => state := s13825; 	--9
	mulfpsclr <= '0';
when s13825 => state := s13826; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13826 => 			--11
	if (mulfprdy = '1') then state := s13827;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13826; end if;
when s13827 => state := s13828; 	--12
	mulfpsclr <= '0';
when s13828 => state := s13829; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13829 => 			--14
	if (addfprdy = '1') then state := s13830;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13829; end if;
when s13830 => state := s13831; 	--15
	addfpsclr <= '0';
when s13831 => state := s13832; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13832 => 			--17
	if (addfprdy = '1') then state := s13833;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13832; end if;
when s13833 => state := s13834; 	--18
	addfpsclr <= '0';
when s13834 => state := s13835; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13835 => 			--20
	if (addfprdy = '1') then state := s13836;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13835; end if;
when s13836 => state := s13837; 	--21
	addfpsclr <= '0';
when s13837 => state := s13838; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (684, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13838 => state := s13839; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1306, 12)); -- offset LSB 1258
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s13839 => state := s13840;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1307, 12)); -- offset MSB 1259
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13840 => state := s13841; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13841 => 			--4
	if (fixed2floatrdy = '1') then state := s13842;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13841; end if;
when s13842 => state := s13843; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13843 => 			--6
	if (mulfprdy = '1') then state := s13844;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13843; end if;
when s13844 => state := s13845; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13845 => 			--8
	if (mulfprdy = '1') then state := s13846;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13845; end if;
when s13846 => state := s13847; 	--9
	mulfpsclr <= '0';
when s13847 => state := s13848; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13848 => 			--11
	if (mulfprdy = '1') then state := s13849;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13848; end if;
when s13849 => state := s13850; 	--12
	mulfpsclr <= '0';
when s13850 => state := s13851; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13851 => 			--14
	if (addfprdy = '1') then state := s13852;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13851; end if;
when s13852 => state := s13853; 	--15
	addfpsclr <= '0';
when s13853 => state := s13854; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13854 => 			--17
	if (addfprdy = '1') then state := s13855;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13854; end if;
when s13855 => state := s13856; 	--18
	addfpsclr <= '0';
when s13856 => state := s13857; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13857 => 			--20
	if (addfprdy = '1') then state := s13858;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13857; end if;
when s13858 => state := s13859; 	--21
	addfpsclr <= '0';
when s13859 => state := s13860; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (685, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13860 => state := s13861; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1308, 12)); -- offset LSB 1260
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s13861 => state := s13862;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1309, 12)); -- offset MSB 1261
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13862 => state := s13863; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13863 => 			--4
	if (fixed2floatrdy = '1') then state := s13864;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13863; end if;
when s13864 => state := s13865; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13865 => 			--6
	if (mulfprdy = '1') then state := s13866;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13865; end if;
when s13866 => state := s13867; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13867 => 			--8
	if (mulfprdy = '1') then state := s13868;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13867; end if;
when s13868 => state := s13869; 	--9
	mulfpsclr <= '0';
when s13869 => state := s13870; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13870 => 			--11
	if (mulfprdy = '1') then state := s13871;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13870; end if;
when s13871 => state := s13872; 	--12
	mulfpsclr <= '0';
when s13872 => state := s13873; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13873 => 			--14
	if (addfprdy = '1') then state := s13874;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13873; end if;
when s13874 => state := s13875; 	--15
	addfpsclr <= '0';
when s13875 => state := s13876; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13876 => 			--17
	if (addfprdy = '1') then state := s13877;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13876; end if;
when s13877 => state := s13878; 	--18
	addfpsclr <= '0';
when s13878 => state := s13879; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13879 => 			--20
	if (addfprdy = '1') then state := s13880;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13879; end if;
when s13880 => state := s13881; 	--21
	addfpsclr <= '0';
when s13881 => state := s13882; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (686, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13882 => state := s13883; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1310, 12)); -- offset LSB 1262
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s13883 => state := s13884;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1311, 12)); -- offset MSB 1263
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13884 => state := s13885; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13885 => 			--4
	if (fixed2floatrdy = '1') then state := s13886;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13885; end if;
when s13886 => state := s13887; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13887 => 			--6
	if (mulfprdy = '1') then state := s13888;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13887; end if;
when s13888 => state := s13889; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13889 => 			--8
	if (mulfprdy = '1') then state := s13890;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13889; end if;
when s13890 => state := s13891; 	--9
	mulfpsclr <= '0';
when s13891 => state := s13892; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13892 => 			--11
	if (mulfprdy = '1') then state := s13893;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13892; end if;
when s13893 => state := s13894; 	--12
	mulfpsclr <= '0';
when s13894 => state := s13895; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13895 => 			--14
	if (addfprdy = '1') then state := s13896;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13895; end if;
when s13896 => state := s13897; 	--15
	addfpsclr <= '0';
when s13897 => state := s13898; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13898 => 			--17
	if (addfprdy = '1') then state := s13899;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13898; end if;
when s13899 => state := s13900; 	--18
	addfpsclr <= '0';
when s13900 => state := s13901; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13901 => 			--20
	if (addfprdy = '1') then state := s13902;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13901; end if;
when s13902 => state := s13903; 	--21
	addfpsclr <= '0';
when s13903 => state := s13904; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (687, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13904 => state := s13905; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1312, 12)); -- offset LSB 1264
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s13905 => state := s13906;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1313, 12)); -- offset MSB 1265
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13906 => state := s13907; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13907 => 			--4
	if (fixed2floatrdy = '1') then state := s13908;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13907; end if;
when s13908 => state := s13909; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13909 => 			--6
	if (mulfprdy = '1') then state := s13910;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13909; end if;
when s13910 => state := s13911; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13911 => 			--8
	if (mulfprdy = '1') then state := s13912;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13911; end if;
when s13912 => state := s13913; 	--9
	mulfpsclr <= '0';
when s13913 => state := s13914; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13914 => 			--11
	if (mulfprdy = '1') then state := s13915;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13914; end if;
when s13915 => state := s13916; 	--12
	mulfpsclr <= '0';
when s13916 => state := s13917; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13917 => 			--14
	if (addfprdy = '1') then state := s13918;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13917; end if;
when s13918 => state := s13919; 	--15
	addfpsclr <= '0';
when s13919 => state := s13920; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13920 => 			--17
	if (addfprdy = '1') then state := s13921;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13920; end if;
when s13921 => state := s13922; 	--18
	addfpsclr <= '0';
when s13922 => state := s13923; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13923 => 			--20
	if (addfprdy = '1') then state := s13924;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13923; end if;
when s13924 => state := s13925; 	--21
	addfpsclr <= '0';
when s13925 => state := s13926; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (688, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13926 => state := s13927; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1314, 12)); -- offset LSB 1266
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s13927 => state := s13928;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1315, 12)); -- offset MSB 1267
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13928 => state := s13929; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13929 => 			--4
	if (fixed2floatrdy = '1') then state := s13930;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13929; end if;
when s13930 => state := s13931; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13931 => 			--6
	if (mulfprdy = '1') then state := s13932;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13931; end if;
when s13932 => state := s13933; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13933 => 			--8
	if (mulfprdy = '1') then state := s13934;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13933; end if;
when s13934 => state := s13935; 	--9
	mulfpsclr <= '0';
when s13935 => state := s13936; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13936 => 			--11
	if (mulfprdy = '1') then state := s13937;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13936; end if;
when s13937 => state := s13938; 	--12
	mulfpsclr <= '0';
when s13938 => state := s13939; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13939 => 			--14
	if (addfprdy = '1') then state := s13940;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13939; end if;
when s13940 => state := s13941; 	--15
	addfpsclr <= '0';
when s13941 => state := s13942; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13942 => 			--17
	if (addfprdy = '1') then state := s13943;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13942; end if;
when s13943 => state := s13944; 	--18
	addfpsclr <= '0';
when s13944 => state := s13945; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13945 => 			--20
	if (addfprdy = '1') then state := s13946;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13945; end if;
when s13946 => state := s13947; 	--21
	addfpsclr <= '0';
when s13947 => state := s13948; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (689, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13948 => state := s13949; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1316, 12)); -- offset LSB 1268
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s13949 => state := s13950;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1317, 12)); -- offset MSB 1269
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13950 => state := s13951; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13951 => 			--4
	if (fixed2floatrdy = '1') then state := s13952;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13951; end if;
when s13952 => state := s13953; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13953 => 			--6
	if (mulfprdy = '1') then state := s13954;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13953; end if;
when s13954 => state := s13955; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13955 => 			--8
	if (mulfprdy = '1') then state := s13956;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13955; end if;
when s13956 => state := s13957; 	--9
	mulfpsclr <= '0';
when s13957 => state := s13958; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13958 => 			--11
	if (mulfprdy = '1') then state := s13959;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13958; end if;
when s13959 => state := s13960; 	--12
	mulfpsclr <= '0';
when s13960 => state := s13961; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13961 => 			--14
	if (addfprdy = '1') then state := s13962;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13961; end if;
when s13962 => state := s13963; 	--15
	addfpsclr <= '0';
when s13963 => state := s13964; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13964 => 			--17
	if (addfprdy = '1') then state := s13965;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13964; end if;
when s13965 => state := s13966; 	--18
	addfpsclr <= '0';
when s13966 => state := s13967; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13967 => 			--20
	if (addfprdy = '1') then state := s13968;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13967; end if;
when s13968 => state := s13969; 	--21
	addfpsclr <= '0';
when s13969 => state := s13970; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (690, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13970 => state := s13971; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1318, 12)); -- offset LSB 1270
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s13971 => state := s13972;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1319, 12)); -- offset MSB 1271
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13972 => state := s13973; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13973 => 			--4
	if (fixed2floatrdy = '1') then state := s13974;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13973; end if;
when s13974 => state := s13975; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13975 => 			--6
	if (mulfprdy = '1') then state := s13976;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13975; end if;
when s13976 => state := s13977; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13977 => 			--8
	if (mulfprdy = '1') then state := s13978;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13977; end if;
when s13978 => state := s13979; 	--9
	mulfpsclr <= '0';
when s13979 => state := s13980; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s13980 => 			--11
	if (mulfprdy = '1') then state := s13981;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13980; end if;
when s13981 => state := s13982; 	--12
	mulfpsclr <= '0';
when s13982 => state := s13983; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s13983 => 			--14
	if (addfprdy = '1') then state := s13984;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13983; end if;
when s13984 => state := s13985; 	--15
	addfpsclr <= '0';
when s13985 => state := s13986; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s13986 => 			--17
	if (addfprdy = '1') then state := s13987;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13986; end if;
when s13987 => state := s13988; 	--18
	addfpsclr <= '0';
when s13988 => state := s13989; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s13989 => 			--20
	if (addfprdy = '1') then state := s13990;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s13989; end if;
when s13990 => state := s13991; 	--21
	addfpsclr <= '0';
when s13991 => state := s13992; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (691, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s13992 => state := s13993; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1320, 12)); -- offset LSB 1272
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s13993 => state := s13994;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1321, 12)); -- offset MSB 1273
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s13994 => state := s13995; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s13995 => 			--4
	if (fixed2floatrdy = '1') then state := s13996;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s13995; end if;
when s13996 => state := s13997; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s13997 => 			--6
	if (mulfprdy = '1') then state := s13998;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13997; end if;
when s13998 => state := s13999; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s13999 => 			--8
	if (mulfprdy = '1') then state := s14000;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s13999; end if;
when s14000 => state := s14001; 	--9
	mulfpsclr <= '0';
when s14001 => state := s14002; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14002 => 			--11
	if (mulfprdy = '1') then state := s14003;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14002; end if;
when s14003 => state := s14004; 	--12
	mulfpsclr <= '0';
when s14004 => state := s14005; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14005 => 			--14
	if (addfprdy = '1') then state := s14006;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14005; end if;
when s14006 => state := s14007; 	--15
	addfpsclr <= '0';
when s14007 => state := s14008; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14008 => 			--17
	if (addfprdy = '1') then state := s14009;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14008; end if;
when s14009 => state := s14010; 	--18
	addfpsclr <= '0';
when s14010 => state := s14011; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14011 => 			--20
	if (addfprdy = '1') then state := s14012;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14011; end if;
when s14012 => state := s14013; 	--21
	addfpsclr <= '0';
when s14013 => state := s14014; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (692, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14014 => state := s14015; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1322, 12)); -- offset LSB 1274
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s14015 => state := s14016;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1323, 12)); -- offset MSB 1275
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14016 => state := s14017; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14017 => 			--4
	if (fixed2floatrdy = '1') then state := s14018;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14017; end if;
when s14018 => state := s14019; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14019 => 			--6
	if (mulfprdy = '1') then state := s14020;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14019; end if;
when s14020 => state := s14021; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14021 => 			--8
	if (mulfprdy = '1') then state := s14022;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14021; end if;
when s14022 => state := s14023; 	--9
	mulfpsclr <= '0';
when s14023 => state := s14024; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14024 => 			--11
	if (mulfprdy = '1') then state := s14025;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14024; end if;
when s14025 => state := s14026; 	--12
	mulfpsclr <= '0';
when s14026 => state := s14027; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14027 => 			--14
	if (addfprdy = '1') then state := s14028;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14027; end if;
when s14028 => state := s14029; 	--15
	addfpsclr <= '0';
when s14029 => state := s14030; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14030 => 			--17
	if (addfprdy = '1') then state := s14031;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14030; end if;
when s14031 => state := s14032; 	--18
	addfpsclr <= '0';
when s14032 => state := s14033; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14033 => 			--20
	if (addfprdy = '1') then state := s14034;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14033; end if;
when s14034 => state := s14035; 	--21
	addfpsclr <= '0';
when s14035 => state := s14036; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (693, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14036 => state := s14037; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1324, 12)); -- offset LSB 1276
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s14037 => state := s14038;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1325, 12)); -- offset MSB 1277
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14038 => state := s14039; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14039 => 			--4
	if (fixed2floatrdy = '1') then state := s14040;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14039; end if;
when s14040 => state := s14041; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14041 => 			--6
	if (mulfprdy = '1') then state := s14042;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14041; end if;
when s14042 => state := s14043; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14043 => 			--8
	if (mulfprdy = '1') then state := s14044;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14043; end if;
when s14044 => state := s14045; 	--9
	mulfpsclr <= '0';
when s14045 => state := s14046; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14046 => 			--11
	if (mulfprdy = '1') then state := s14047;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14046; end if;
when s14047 => state := s14048; 	--12
	mulfpsclr <= '0';
when s14048 => state := s14049; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14049 => 			--14
	if (addfprdy = '1') then state := s14050;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14049; end if;
when s14050 => state := s14051; 	--15
	addfpsclr <= '0';
when s14051 => state := s14052; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14052 => 			--17
	if (addfprdy = '1') then state := s14053;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14052; end if;
when s14053 => state := s14054; 	--18
	addfpsclr <= '0';
when s14054 => state := s14055; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14055 => 			--20
	if (addfprdy = '1') then state := s14056;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14055; end if;
when s14056 => state := s14057; 	--21
	addfpsclr <= '0';
when s14057 => state := s14058; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (694, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14058 => state := s14059; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1326, 12)); -- offset LSB 1278
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s14059 => state := s14060;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1327, 12)); -- offset MSB 1279
	addra <= std_logic_vector (to_unsigned (19, 10)); -- OCCrowI 19
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14060 => state := s14061; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14061 => 			--4
	if (fixed2floatrdy = '1') then state := s14062;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14061; end if;
when s14062 => state := s14063; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14063 => 			--6
	if (mulfprdy = '1') then state := s14064;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14063; end if;
when s14064 => state := s14065; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14065 => 			--8
	if (mulfprdy = '1') then state := s14066;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14065; end if;
when s14066 => state := s14067; 	--9
	mulfpsclr <= '0';
when s14067 => state := s14068; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14068 => 			--11
	if (mulfprdy = '1') then state := s14069;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14068; end if;
when s14069 => state := s14070; 	--12
	mulfpsclr <= '0';
when s14070 => state := s14071; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14071 => 			--14
	if (addfprdy = '1') then state := s14072;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14071; end if;
when s14072 => state := s14073; 	--15
	addfpsclr <= '0';
when s14073 => state := s14074; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14074 => 			--17
	if (addfprdy = '1') then state := s14075;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14074; end if;
when s14075 => state := s14076; 	--18
	addfpsclr <= '0';
when s14076 => state := s14077; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14077 => 			--20
	if (addfprdy = '1') then state := s14078;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14077; end if;
when s14078 => state := s14079; 	--21
	addfpsclr <= '0';
when s14079 => state := s14080; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (695, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14080 => state := s14081; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1328, 12)); -- offset LSB 1280
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s14081 => state := s14082;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1329, 12)); -- offset MSB 1281
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14082 => state := s14083; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14083 => 			--4
	if (fixed2floatrdy = '1') then state := s14084;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14083; end if;
when s14084 => state := s14085; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14085 => 			--6
	if (mulfprdy = '1') then state := s14086;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14085; end if;
when s14086 => state := s14087; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14087 => 			--8
	if (mulfprdy = '1') then state := s14088;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14087; end if;
when s14088 => state := s14089; 	--9
	mulfpsclr <= '0';
when s14089 => state := s14090; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14090 => 			--11
	if (mulfprdy = '1') then state := s14091;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14090; end if;
when s14091 => state := s14092; 	--12
	mulfpsclr <= '0';
when s14092 => state := s14093; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14093 => 			--14
	if (addfprdy = '1') then state := s14094;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14093; end if;
when s14094 => state := s14095; 	--15
	addfpsclr <= '0';
when s14095 => state := s14096; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14096 => 			--17
	if (addfprdy = '1') then state := s14097;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14096; end if;
when s14097 => state := s14098; 	--18
	addfpsclr <= '0';
when s14098 => state := s14099; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14099 => 			--20
	if (addfprdy = '1') then state := s14100;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14099; end if;
when s14100 => state := s14101; 	--21
	addfpsclr <= '0';
when s14101 => state := s14102; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (696, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14102 => state := s14103; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1330, 12)); -- offset LSB 1282
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s14103 => state := s14104;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1331, 12)); -- offset MSB 1283
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14104 => state := s14105; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14105 => 			--4
	if (fixed2floatrdy = '1') then state := s14106;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14105; end if;
when s14106 => state := s14107; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14107 => 			--6
	if (mulfprdy = '1') then state := s14108;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14107; end if;
when s14108 => state := s14109; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14109 => 			--8
	if (mulfprdy = '1') then state := s14110;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14109; end if;
when s14110 => state := s14111; 	--9
	mulfpsclr <= '0';
when s14111 => state := s14112; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14112 => 			--11
	if (mulfprdy = '1') then state := s14113;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14112; end if;
when s14113 => state := s14114; 	--12
	mulfpsclr <= '0';
when s14114 => state := s14115; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14115 => 			--14
	if (addfprdy = '1') then state := s14116;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14115; end if;
when s14116 => state := s14117; 	--15
	addfpsclr <= '0';
when s14117 => state := s14118; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14118 => 			--17
	if (addfprdy = '1') then state := s14119;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14118; end if;
when s14119 => state := s14120; 	--18
	addfpsclr <= '0';
when s14120 => state := s14121; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14121 => 			--20
	if (addfprdy = '1') then state := s14122;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14121; end if;
when s14122 => state := s14123; 	--21
	addfpsclr <= '0';
when s14123 => state := s14124; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (697, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14124 => state := s14125; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1332, 12)); -- offset LSB 1284
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s14125 => state := s14126;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1333, 12)); -- offset MSB 1285
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14126 => state := s14127; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14127 => 			--4
	if (fixed2floatrdy = '1') then state := s14128;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14127; end if;
when s14128 => state := s14129; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14129 => 			--6
	if (mulfprdy = '1') then state := s14130;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14129; end if;
when s14130 => state := s14131; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14131 => 			--8
	if (mulfprdy = '1') then state := s14132;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14131; end if;
when s14132 => state := s14133; 	--9
	mulfpsclr <= '0';
when s14133 => state := s14134; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14134 => 			--11
	if (mulfprdy = '1') then state := s14135;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14134; end if;
when s14135 => state := s14136; 	--12
	mulfpsclr <= '0';
when s14136 => state := s14137; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14137 => 			--14
	if (addfprdy = '1') then state := s14138;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14137; end if;
when s14138 => state := s14139; 	--15
	addfpsclr <= '0';
when s14139 => state := s14140; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14140 => 			--17
	if (addfprdy = '1') then state := s14141;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14140; end if;
when s14141 => state := s14142; 	--18
	addfpsclr <= '0';
when s14142 => state := s14143; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14143 => 			--20
	if (addfprdy = '1') then state := s14144;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14143; end if;
when s14144 => state := s14145; 	--21
	addfpsclr <= '0';
when s14145 => state := s14146; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (698, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14146 => state := s14147; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1334, 12)); -- offset LSB 1286
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s14147 => state := s14148;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1335, 12)); -- offset MSB 1287
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14148 => state := s14149; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14149 => 			--4
	if (fixed2floatrdy = '1') then state := s14150;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14149; end if;
when s14150 => state := s14151; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14151 => 			--6
	if (mulfprdy = '1') then state := s14152;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14151; end if;
when s14152 => state := s14153; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14153 => 			--8
	if (mulfprdy = '1') then state := s14154;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14153; end if;
when s14154 => state := s14155; 	--9
	mulfpsclr <= '0';
when s14155 => state := s14156; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14156 => 			--11
	if (mulfprdy = '1') then state := s14157;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14156; end if;
when s14157 => state := s14158; 	--12
	mulfpsclr <= '0';
when s14158 => state := s14159; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14159 => 			--14
	if (addfprdy = '1') then state := s14160;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14159; end if;
when s14160 => state := s14161; 	--15
	addfpsclr <= '0';
when s14161 => state := s14162; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14162 => 			--17
	if (addfprdy = '1') then state := s14163;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14162; end if;
when s14163 => state := s14164; 	--18
	addfpsclr <= '0';
when s14164 => state := s14165; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14165 => 			--20
	if (addfprdy = '1') then state := s14166;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14165; end if;
when s14166 => state := s14167; 	--21
	addfpsclr <= '0';
when s14167 => state := s14168; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (699, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14168 => state := s14169; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1336, 12)); -- offset LSB 1288
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s14169 => state := s14170;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1337, 12)); -- offset MSB 1289
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14170 => state := s14171; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14171 => 			--4
	if (fixed2floatrdy = '1') then state := s14172;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14171; end if;
when s14172 => state := s14173; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14173 => 			--6
	if (mulfprdy = '1') then state := s14174;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14173; end if;
when s14174 => state := s14175; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14175 => 			--8
	if (mulfprdy = '1') then state := s14176;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14175; end if;
when s14176 => state := s14177; 	--9
	mulfpsclr <= '0';
when s14177 => state := s14178; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14178 => 			--11
	if (mulfprdy = '1') then state := s14179;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14178; end if;
when s14179 => state := s14180; 	--12
	mulfpsclr <= '0';
when s14180 => state := s14181; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14181 => 			--14
	if (addfprdy = '1') then state := s14182;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14181; end if;
when s14182 => state := s14183; 	--15
	addfpsclr <= '0';
when s14183 => state := s14184; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14184 => 			--17
	if (addfprdy = '1') then state := s14185;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14184; end if;
when s14185 => state := s14186; 	--18
	addfpsclr <= '0';
when s14186 => state := s14187; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14187 => 			--20
	if (addfprdy = '1') then state := s14188;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14187; end if;
when s14188 => state := s14189; 	--21
	addfpsclr <= '0';
when s14189 => state := s14190; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (700, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14190 => state := s14191; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1338, 12)); -- offset LSB 1290
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s14191 => state := s14192;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1339, 12)); -- offset MSB 1291
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14192 => state := s14193; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14193 => 			--4
	if (fixed2floatrdy = '1') then state := s14194;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14193; end if;
when s14194 => state := s14195; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14195 => 			--6
	if (mulfprdy = '1') then state := s14196;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14195; end if;
when s14196 => state := s14197; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14197 => 			--8
	if (mulfprdy = '1') then state := s14198;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14197; end if;
when s14198 => state := s14199; 	--9
	mulfpsclr <= '0';
when s14199 => state := s14200; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14200 => 			--11
	if (mulfprdy = '1') then state := s14201;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14200; end if;
when s14201 => state := s14202; 	--12
	mulfpsclr <= '0';
when s14202 => state := s14203; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14203 => 			--14
	if (addfprdy = '1') then state := s14204;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14203; end if;
when s14204 => state := s14205; 	--15
	addfpsclr <= '0';
when s14205 => state := s14206; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14206 => 			--17
	if (addfprdy = '1') then state := s14207;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14206; end if;
when s14207 => state := s14208; 	--18
	addfpsclr <= '0';
when s14208 => state := s14209; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14209 => 			--20
	if (addfprdy = '1') then state := s14210;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14209; end if;
when s14210 => state := s14211; 	--21
	addfpsclr <= '0';
when s14211 => state := s14212; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (701, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14212 => state := s14213; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1340, 12)); -- offset LSB 1292
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s14213 => state := s14214;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1341, 12)); -- offset MSB 1293
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14214 => state := s14215; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14215 => 			--4
	if (fixed2floatrdy = '1') then state := s14216;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14215; end if;
when s14216 => state := s14217; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14217 => 			--6
	if (mulfprdy = '1') then state := s14218;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14217; end if;
when s14218 => state := s14219; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14219 => 			--8
	if (mulfprdy = '1') then state := s14220;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14219; end if;
when s14220 => state := s14221; 	--9
	mulfpsclr <= '0';
when s14221 => state := s14222; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14222 => 			--11
	if (mulfprdy = '1') then state := s14223;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14222; end if;
when s14223 => state := s14224; 	--12
	mulfpsclr <= '0';
when s14224 => state := s14225; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14225 => 			--14
	if (addfprdy = '1') then state := s14226;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14225; end if;
when s14226 => state := s14227; 	--15
	addfpsclr <= '0';
when s14227 => state := s14228; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14228 => 			--17
	if (addfprdy = '1') then state := s14229;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14228; end if;
when s14229 => state := s14230; 	--18
	addfpsclr <= '0';
when s14230 => state := s14231; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14231 => 			--20
	if (addfprdy = '1') then state := s14232;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14231; end if;
when s14232 => state := s14233; 	--21
	addfpsclr <= '0';
when s14233 => state := s14234; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (702, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14234 => state := s14235; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1342, 12)); -- offset LSB 1294
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s14235 => state := s14236;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1343, 12)); -- offset MSB 1295
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14236 => state := s14237; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14237 => 			--4
	if (fixed2floatrdy = '1') then state := s14238;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14237; end if;
when s14238 => state := s14239; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14239 => 			--6
	if (mulfprdy = '1') then state := s14240;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14239; end if;
when s14240 => state := s14241; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14241 => 			--8
	if (mulfprdy = '1') then state := s14242;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14241; end if;
when s14242 => state := s14243; 	--9
	mulfpsclr <= '0';
when s14243 => state := s14244; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14244 => 			--11
	if (mulfprdy = '1') then state := s14245;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14244; end if;
when s14245 => state := s14246; 	--12
	mulfpsclr <= '0';
when s14246 => state := s14247; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14247 => 			--14
	if (addfprdy = '1') then state := s14248;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14247; end if;
when s14248 => state := s14249; 	--15
	addfpsclr <= '0';
when s14249 => state := s14250; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14250 => 			--17
	if (addfprdy = '1') then state := s14251;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14250; end if;
when s14251 => state := s14252; 	--18
	addfpsclr <= '0';
when s14252 => state := s14253; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14253 => 			--20
	if (addfprdy = '1') then state := s14254;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14253; end if;
when s14254 => state := s14255; 	--21
	addfpsclr <= '0';
when s14255 => state := s14256; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (703, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14256 => state := s14257; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1344, 12)); -- offset LSB 1296
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s14257 => state := s14258;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1345, 12)); -- offset MSB 1297
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14258 => state := s14259; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14259 => 			--4
	if (fixed2floatrdy = '1') then state := s14260;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14259; end if;
when s14260 => state := s14261; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14261 => 			--6
	if (mulfprdy = '1') then state := s14262;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14261; end if;
when s14262 => state := s14263; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14263 => 			--8
	if (mulfprdy = '1') then state := s14264;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14263; end if;
when s14264 => state := s14265; 	--9
	mulfpsclr <= '0';
when s14265 => state := s14266; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14266 => 			--11
	if (mulfprdy = '1') then state := s14267;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14266; end if;
when s14267 => state := s14268; 	--12
	mulfpsclr <= '0';
when s14268 => state := s14269; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14269 => 			--14
	if (addfprdy = '1') then state := s14270;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14269; end if;
when s14270 => state := s14271; 	--15
	addfpsclr <= '0';
when s14271 => state := s14272; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14272 => 			--17
	if (addfprdy = '1') then state := s14273;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14272; end if;
when s14273 => state := s14274; 	--18
	addfpsclr <= '0';
when s14274 => state := s14275; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14275 => 			--20
	if (addfprdy = '1') then state := s14276;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14275; end if;
when s14276 => state := s14277; 	--21
	addfpsclr <= '0';
when s14277 => state := s14278; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (704, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14278 => state := s14279; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1346, 12)); -- offset LSB 1298
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s14279 => state := s14280;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1347, 12)); -- offset MSB 1299
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14280 => state := s14281; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14281 => 			--4
	if (fixed2floatrdy = '1') then state := s14282;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14281; end if;
when s14282 => state := s14283; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14283 => 			--6
	if (mulfprdy = '1') then state := s14284;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14283; end if;
when s14284 => state := s14285; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14285 => 			--8
	if (mulfprdy = '1') then state := s14286;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14285; end if;
when s14286 => state := s14287; 	--9
	mulfpsclr <= '0';
when s14287 => state := s14288; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14288 => 			--11
	if (mulfprdy = '1') then state := s14289;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14288; end if;
when s14289 => state := s14290; 	--12
	mulfpsclr <= '0';
when s14290 => state := s14291; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14291 => 			--14
	if (addfprdy = '1') then state := s14292;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14291; end if;
when s14292 => state := s14293; 	--15
	addfpsclr <= '0';
when s14293 => state := s14294; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14294 => 			--17
	if (addfprdy = '1') then state := s14295;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14294; end if;
when s14295 => state := s14296; 	--18
	addfpsclr <= '0';
when s14296 => state := s14297; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14297 => 			--20
	if (addfprdy = '1') then state := s14298;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14297; end if;
when s14298 => state := s14299; 	--21
	addfpsclr <= '0';
when s14299 => state := s14300; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (705, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14300 => state := s14301; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1348, 12)); -- offset LSB 1300
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s14301 => state := s14302;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1349, 12)); -- offset MSB 1301
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14302 => state := s14303; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14303 => 			--4
	if (fixed2floatrdy = '1') then state := s14304;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14303; end if;
when s14304 => state := s14305; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14305 => 			--6
	if (mulfprdy = '1') then state := s14306;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14305; end if;
when s14306 => state := s14307; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14307 => 			--8
	if (mulfprdy = '1') then state := s14308;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14307; end if;
when s14308 => state := s14309; 	--9
	mulfpsclr <= '0';
when s14309 => state := s14310; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14310 => 			--11
	if (mulfprdy = '1') then state := s14311;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14310; end if;
when s14311 => state := s14312; 	--12
	mulfpsclr <= '0';
when s14312 => state := s14313; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14313 => 			--14
	if (addfprdy = '1') then state := s14314;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14313; end if;
when s14314 => state := s14315; 	--15
	addfpsclr <= '0';
when s14315 => state := s14316; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14316 => 			--17
	if (addfprdy = '1') then state := s14317;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14316; end if;
when s14317 => state := s14318; 	--18
	addfpsclr <= '0';
when s14318 => state := s14319; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14319 => 			--20
	if (addfprdy = '1') then state := s14320;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14319; end if;
when s14320 => state := s14321; 	--21
	addfpsclr <= '0';
when s14321 => state := s14322; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (706, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14322 => state := s14323; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1350, 12)); -- offset LSB 1302
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s14323 => state := s14324;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1351, 12)); -- offset MSB 1303
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14324 => state := s14325; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14325 => 			--4
	if (fixed2floatrdy = '1') then state := s14326;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14325; end if;
when s14326 => state := s14327; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14327 => 			--6
	if (mulfprdy = '1') then state := s14328;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14327; end if;
when s14328 => state := s14329; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14329 => 			--8
	if (mulfprdy = '1') then state := s14330;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14329; end if;
when s14330 => state := s14331; 	--9
	mulfpsclr <= '0';
when s14331 => state := s14332; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14332 => 			--11
	if (mulfprdy = '1') then state := s14333;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14332; end if;
when s14333 => state := s14334; 	--12
	mulfpsclr <= '0';
when s14334 => state := s14335; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14335 => 			--14
	if (addfprdy = '1') then state := s14336;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14335; end if;
when s14336 => state := s14337; 	--15
	addfpsclr <= '0';
when s14337 => state := s14338; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14338 => 			--17
	if (addfprdy = '1') then state := s14339;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14338; end if;
when s14339 => state := s14340; 	--18
	addfpsclr <= '0';
when s14340 => state := s14341; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14341 => 			--20
	if (addfprdy = '1') then state := s14342;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14341; end if;
when s14342 => state := s14343; 	--21
	addfpsclr <= '0';
when s14343 => state := s14344; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (707, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14344 => state := s14345; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1352, 12)); -- offset LSB 1304
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s14345 => state := s14346;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1353, 12)); -- offset MSB 1305
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14346 => state := s14347; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14347 => 			--4
	if (fixed2floatrdy = '1') then state := s14348;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14347; end if;
when s14348 => state := s14349; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14349 => 			--6
	if (mulfprdy = '1') then state := s14350;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14349; end if;
when s14350 => state := s14351; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14351 => 			--8
	if (mulfprdy = '1') then state := s14352;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14351; end if;
when s14352 => state := s14353; 	--9
	mulfpsclr <= '0';
when s14353 => state := s14354; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14354 => 			--11
	if (mulfprdy = '1') then state := s14355;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14354; end if;
when s14355 => state := s14356; 	--12
	mulfpsclr <= '0';
when s14356 => state := s14357; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14357 => 			--14
	if (addfprdy = '1') then state := s14358;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14357; end if;
when s14358 => state := s14359; 	--15
	addfpsclr <= '0';
when s14359 => state := s14360; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14360 => 			--17
	if (addfprdy = '1') then state := s14361;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14360; end if;
when s14361 => state := s14362; 	--18
	addfpsclr <= '0';
when s14362 => state := s14363; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14363 => 			--20
	if (addfprdy = '1') then state := s14364;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14363; end if;
when s14364 => state := s14365; 	--21
	addfpsclr <= '0';
when s14365 => state := s14366; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (708, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14366 => state := s14367; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1354, 12)); -- offset LSB 1306
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s14367 => state := s14368;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1355, 12)); -- offset MSB 1307
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14368 => state := s14369; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14369 => 			--4
	if (fixed2floatrdy = '1') then state := s14370;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14369; end if;
when s14370 => state := s14371; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14371 => 			--6
	if (mulfprdy = '1') then state := s14372;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14371; end if;
when s14372 => state := s14373; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14373 => 			--8
	if (mulfprdy = '1') then state := s14374;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14373; end if;
when s14374 => state := s14375; 	--9
	mulfpsclr <= '0';
when s14375 => state := s14376; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14376 => 			--11
	if (mulfprdy = '1') then state := s14377;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14376; end if;
when s14377 => state := s14378; 	--12
	mulfpsclr <= '0';
when s14378 => state := s14379; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14379 => 			--14
	if (addfprdy = '1') then state := s14380;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14379; end if;
when s14380 => state := s14381; 	--15
	addfpsclr <= '0';
when s14381 => state := s14382; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14382 => 			--17
	if (addfprdy = '1') then state := s14383;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14382; end if;
when s14383 => state := s14384; 	--18
	addfpsclr <= '0';
when s14384 => state := s14385; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14385 => 			--20
	if (addfprdy = '1') then state := s14386;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14385; end if;
when s14386 => state := s14387; 	--21
	addfpsclr <= '0';
when s14387 => state := s14388; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (709, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14388 => state := s14389; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1356, 12)); -- offset LSB 1308
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s14389 => state := s14390;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1357, 12)); -- offset MSB 1309
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14390 => state := s14391; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14391 => 			--4
	if (fixed2floatrdy = '1') then state := s14392;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14391; end if;
when s14392 => state := s14393; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14393 => 			--6
	if (mulfprdy = '1') then state := s14394;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14393; end if;
when s14394 => state := s14395; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14395 => 			--8
	if (mulfprdy = '1') then state := s14396;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14395; end if;
when s14396 => state := s14397; 	--9
	mulfpsclr <= '0';
when s14397 => state := s14398; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14398 => 			--11
	if (mulfprdy = '1') then state := s14399;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14398; end if;
when s14399 => state := s14400; 	--12
	mulfpsclr <= '0';
when s14400 => state := s14401; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14401 => 			--14
	if (addfprdy = '1') then state := s14402;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14401; end if;
when s14402 => state := s14403; 	--15
	addfpsclr <= '0';
when s14403 => state := s14404; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14404 => 			--17
	if (addfprdy = '1') then state := s14405;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14404; end if;
when s14405 => state := s14406; 	--18
	addfpsclr <= '0';
when s14406 => state := s14407; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14407 => 			--20
	if (addfprdy = '1') then state := s14408;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14407; end if;
when s14408 => state := s14409; 	--21
	addfpsclr <= '0';
when s14409 => state := s14410; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (710, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14410 => state := s14411; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1358, 12)); -- offset LSB 1310
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s14411 => state := s14412;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1359, 12)); -- offset MSB 1311
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14412 => state := s14413; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14413 => 			--4
	if (fixed2floatrdy = '1') then state := s14414;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14413; end if;
when s14414 => state := s14415; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14415 => 			--6
	if (mulfprdy = '1') then state := s14416;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14415; end if;
when s14416 => state := s14417; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14417 => 			--8
	if (mulfprdy = '1') then state := s14418;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14417; end if;
when s14418 => state := s14419; 	--9
	mulfpsclr <= '0';
when s14419 => state := s14420; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14420 => 			--11
	if (mulfprdy = '1') then state := s14421;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14420; end if;
when s14421 => state := s14422; 	--12
	mulfpsclr <= '0';
when s14422 => state := s14423; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14423 => 			--14
	if (addfprdy = '1') then state := s14424;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14423; end if;
when s14424 => state := s14425; 	--15
	addfpsclr <= '0';
when s14425 => state := s14426; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14426 => 			--17
	if (addfprdy = '1') then state := s14427;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14426; end if;
when s14427 => state := s14428; 	--18
	addfpsclr <= '0';
when s14428 => state := s14429; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14429 => 			--20
	if (addfprdy = '1') then state := s14430;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14429; end if;
when s14430 => state := s14431; 	--21
	addfpsclr <= '0';
when s14431 => state := s14432; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (711, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14432 => state := s14433; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1360, 12)); -- offset LSB 1312
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s14433 => state := s14434;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1361, 12)); -- offset MSB 1313
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14434 => state := s14435; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14435 => 			--4
	if (fixed2floatrdy = '1') then state := s14436;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14435; end if;
when s14436 => state := s14437; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14437 => 			--6
	if (mulfprdy = '1') then state := s14438;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14437; end if;
when s14438 => state := s14439; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14439 => 			--8
	if (mulfprdy = '1') then state := s14440;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14439; end if;
when s14440 => state := s14441; 	--9
	mulfpsclr <= '0';
when s14441 => state := s14442; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14442 => 			--11
	if (mulfprdy = '1') then state := s14443;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14442; end if;
when s14443 => state := s14444; 	--12
	mulfpsclr <= '0';
when s14444 => state := s14445; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14445 => 			--14
	if (addfprdy = '1') then state := s14446;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14445; end if;
when s14446 => state := s14447; 	--15
	addfpsclr <= '0';
when s14447 => state := s14448; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14448 => 			--17
	if (addfprdy = '1') then state := s14449;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14448; end if;
when s14449 => state := s14450; 	--18
	addfpsclr <= '0';
when s14450 => state := s14451; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14451 => 			--20
	if (addfprdy = '1') then state := s14452;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14451; end if;
when s14452 => state := s14453; 	--21
	addfpsclr <= '0';
when s14453 => state := s14454; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (712, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14454 => state := s14455; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1362, 12)); -- offset LSB 1314
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s14455 => state := s14456;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1363, 12)); -- offset MSB 1315
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14456 => state := s14457; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14457 => 			--4
	if (fixed2floatrdy = '1') then state := s14458;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14457; end if;
when s14458 => state := s14459; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14459 => 			--6
	if (mulfprdy = '1') then state := s14460;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14459; end if;
when s14460 => state := s14461; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14461 => 			--8
	if (mulfprdy = '1') then state := s14462;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14461; end if;
when s14462 => state := s14463; 	--9
	mulfpsclr <= '0';
when s14463 => state := s14464; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14464 => 			--11
	if (mulfprdy = '1') then state := s14465;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14464; end if;
when s14465 => state := s14466; 	--12
	mulfpsclr <= '0';
when s14466 => state := s14467; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14467 => 			--14
	if (addfprdy = '1') then state := s14468;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14467; end if;
when s14468 => state := s14469; 	--15
	addfpsclr <= '0';
when s14469 => state := s14470; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14470 => 			--17
	if (addfprdy = '1') then state := s14471;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14470; end if;
when s14471 => state := s14472; 	--18
	addfpsclr <= '0';
when s14472 => state := s14473; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14473 => 			--20
	if (addfprdy = '1') then state := s14474;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14473; end if;
when s14474 => state := s14475; 	--21
	addfpsclr <= '0';
when s14475 => state := s14476; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (713, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14476 => state := s14477; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1364, 12)); -- offset LSB 1316
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s14477 => state := s14478;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1365, 12)); -- offset MSB 1317
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14478 => state := s14479; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14479 => 			--4
	if (fixed2floatrdy = '1') then state := s14480;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14479; end if;
when s14480 => state := s14481; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14481 => 			--6
	if (mulfprdy = '1') then state := s14482;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14481; end if;
when s14482 => state := s14483; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14483 => 			--8
	if (mulfprdy = '1') then state := s14484;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14483; end if;
when s14484 => state := s14485; 	--9
	mulfpsclr <= '0';
when s14485 => state := s14486; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14486 => 			--11
	if (mulfprdy = '1') then state := s14487;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14486; end if;
when s14487 => state := s14488; 	--12
	mulfpsclr <= '0';
when s14488 => state := s14489; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14489 => 			--14
	if (addfprdy = '1') then state := s14490;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14489; end if;
when s14490 => state := s14491; 	--15
	addfpsclr <= '0';
when s14491 => state := s14492; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14492 => 			--17
	if (addfprdy = '1') then state := s14493;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14492; end if;
when s14493 => state := s14494; 	--18
	addfpsclr <= '0';
when s14494 => state := s14495; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14495 => 			--20
	if (addfprdy = '1') then state := s14496;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14495; end if;
when s14496 => state := s14497; 	--21
	addfpsclr <= '0';
when s14497 => state := s14498; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (714, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14498 => state := s14499; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1366, 12)); -- offset LSB 1318
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s14499 => state := s14500;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1367, 12)); -- offset MSB 1319
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14500 => state := s14501; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14501 => 			--4
	if (fixed2floatrdy = '1') then state := s14502;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14501; end if;
when s14502 => state := s14503; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14503 => 			--6
	if (mulfprdy = '1') then state := s14504;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14503; end if;
when s14504 => state := s14505; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14505 => 			--8
	if (mulfprdy = '1') then state := s14506;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14505; end if;
when s14506 => state := s14507; 	--9
	mulfpsclr <= '0';
when s14507 => state := s14508; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14508 => 			--11
	if (mulfprdy = '1') then state := s14509;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14508; end if;
when s14509 => state := s14510; 	--12
	mulfpsclr <= '0';
when s14510 => state := s14511; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14511 => 			--14
	if (addfprdy = '1') then state := s14512;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14511; end if;
when s14512 => state := s14513; 	--15
	addfpsclr <= '0';
when s14513 => state := s14514; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14514 => 			--17
	if (addfprdy = '1') then state := s14515;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14514; end if;
when s14515 => state := s14516; 	--18
	addfpsclr <= '0';
when s14516 => state := s14517; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14517 => 			--20
	if (addfprdy = '1') then state := s14518;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14517; end if;
when s14518 => state := s14519; 	--21
	addfpsclr <= '0';
when s14519 => state := s14520; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (715, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14520 => state := s14521; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1368, 12)); -- offset LSB 1320
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s14521 => state := s14522;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1369, 12)); -- offset MSB 1321
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14522 => state := s14523; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14523 => 			--4
	if (fixed2floatrdy = '1') then state := s14524;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14523; end if;
when s14524 => state := s14525; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14525 => 			--6
	if (mulfprdy = '1') then state := s14526;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14525; end if;
when s14526 => state := s14527; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14527 => 			--8
	if (mulfprdy = '1') then state := s14528;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14527; end if;
when s14528 => state := s14529; 	--9
	mulfpsclr <= '0';
when s14529 => state := s14530; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14530 => 			--11
	if (mulfprdy = '1') then state := s14531;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14530; end if;
when s14531 => state := s14532; 	--12
	mulfpsclr <= '0';
when s14532 => state := s14533; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14533 => 			--14
	if (addfprdy = '1') then state := s14534;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14533; end if;
when s14534 => state := s14535; 	--15
	addfpsclr <= '0';
when s14535 => state := s14536; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14536 => 			--17
	if (addfprdy = '1') then state := s14537;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14536; end if;
when s14537 => state := s14538; 	--18
	addfpsclr <= '0';
when s14538 => state := s14539; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14539 => 			--20
	if (addfprdy = '1') then state := s14540;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14539; end if;
when s14540 => state := s14541; 	--21
	addfpsclr <= '0';
when s14541 => state := s14542; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (716, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14542 => state := s14543; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1370, 12)); -- offset LSB 1322
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s14543 => state := s14544;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1371, 12)); -- offset MSB 1323
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14544 => state := s14545; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14545 => 			--4
	if (fixed2floatrdy = '1') then state := s14546;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14545; end if;
when s14546 => state := s14547; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14547 => 			--6
	if (mulfprdy = '1') then state := s14548;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14547; end if;
when s14548 => state := s14549; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14549 => 			--8
	if (mulfprdy = '1') then state := s14550;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14549; end if;
when s14550 => state := s14551; 	--9
	mulfpsclr <= '0';
when s14551 => state := s14552; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14552 => 			--11
	if (mulfprdy = '1') then state := s14553;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14552; end if;
when s14553 => state := s14554; 	--12
	mulfpsclr <= '0';
when s14554 => state := s14555; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14555 => 			--14
	if (addfprdy = '1') then state := s14556;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14555; end if;
when s14556 => state := s14557; 	--15
	addfpsclr <= '0';
when s14557 => state := s14558; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14558 => 			--17
	if (addfprdy = '1') then state := s14559;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14558; end if;
when s14559 => state := s14560; 	--18
	addfpsclr <= '0';
when s14560 => state := s14561; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14561 => 			--20
	if (addfprdy = '1') then state := s14562;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14561; end if;
when s14562 => state := s14563; 	--21
	addfpsclr <= '0';
when s14563 => state := s14564; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (717, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14564 => state := s14565; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1372, 12)); -- offset LSB 1324
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s14565 => state := s14566;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1373, 12)); -- offset MSB 1325
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14566 => state := s14567; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14567 => 			--4
	if (fixed2floatrdy = '1') then state := s14568;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14567; end if;
when s14568 => state := s14569; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14569 => 			--6
	if (mulfprdy = '1') then state := s14570;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14569; end if;
when s14570 => state := s14571; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14571 => 			--8
	if (mulfprdy = '1') then state := s14572;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14571; end if;
when s14572 => state := s14573; 	--9
	mulfpsclr <= '0';
when s14573 => state := s14574; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14574 => 			--11
	if (mulfprdy = '1') then state := s14575;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14574; end if;
when s14575 => state := s14576; 	--12
	mulfpsclr <= '0';
when s14576 => state := s14577; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14577 => 			--14
	if (addfprdy = '1') then state := s14578;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14577; end if;
when s14578 => state := s14579; 	--15
	addfpsclr <= '0';
when s14579 => state := s14580; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14580 => 			--17
	if (addfprdy = '1') then state := s14581;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14580; end if;
when s14581 => state := s14582; 	--18
	addfpsclr <= '0';
when s14582 => state := s14583; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14583 => 			--20
	if (addfprdy = '1') then state := s14584;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14583; end if;
when s14584 => state := s14585; 	--21
	addfpsclr <= '0';
when s14585 => state := s14586; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (718, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14586 => state := s14587; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1374, 12)); -- offset LSB 1326
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s14587 => state := s14588;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1375, 12)); -- offset MSB 1327
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14588 => state := s14589; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14589 => 			--4
	if (fixed2floatrdy = '1') then state := s14590;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14589; end if;
when s14590 => state := s14591; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14591 => 			--6
	if (mulfprdy = '1') then state := s14592;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14591; end if;
when s14592 => state := s14593; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14593 => 			--8
	if (mulfprdy = '1') then state := s14594;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14593; end if;
when s14594 => state := s14595; 	--9
	mulfpsclr <= '0';
when s14595 => state := s14596; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14596 => 			--11
	if (mulfprdy = '1') then state := s14597;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14596; end if;
when s14597 => state := s14598; 	--12
	mulfpsclr <= '0';
when s14598 => state := s14599; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14599 => 			--14
	if (addfprdy = '1') then state := s14600;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14599; end if;
when s14600 => state := s14601; 	--15
	addfpsclr <= '0';
when s14601 => state := s14602; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14602 => 			--17
	if (addfprdy = '1') then state := s14603;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14602; end if;
when s14603 => state := s14604; 	--18
	addfpsclr <= '0';
when s14604 => state := s14605; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14605 => 			--20
	if (addfprdy = '1') then state := s14606;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14605; end if;
when s14606 => state := s14607; 	--21
	addfpsclr <= '0';
when s14607 => state := s14608; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (719, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14608 => state := s14609; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1376, 12)); -- offset LSB 1328
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s14609 => state := s14610;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1377, 12)); -- offset MSB 1329
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14610 => state := s14611; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14611 => 			--4
	if (fixed2floatrdy = '1') then state := s14612;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14611; end if;
when s14612 => state := s14613; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14613 => 			--6
	if (mulfprdy = '1') then state := s14614;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14613; end if;
when s14614 => state := s14615; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14615 => 			--8
	if (mulfprdy = '1') then state := s14616;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14615; end if;
when s14616 => state := s14617; 	--9
	mulfpsclr <= '0';
when s14617 => state := s14618; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14618 => 			--11
	if (mulfprdy = '1') then state := s14619;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14618; end if;
when s14619 => state := s14620; 	--12
	mulfpsclr <= '0';
when s14620 => state := s14621; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14621 => 			--14
	if (addfprdy = '1') then state := s14622;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14621; end if;
when s14622 => state := s14623; 	--15
	addfpsclr <= '0';
when s14623 => state := s14624; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14624 => 			--17
	if (addfprdy = '1') then state := s14625;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14624; end if;
when s14625 => state := s14626; 	--18
	addfpsclr <= '0';
when s14626 => state := s14627; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14627 => 			--20
	if (addfprdy = '1') then state := s14628;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14627; end if;
when s14628 => state := s14629; 	--21
	addfpsclr <= '0';
when s14629 => state := s14630; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (720, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14630 => state := s14631; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1378, 12)); -- offset LSB 1330
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s14631 => state := s14632;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1379, 12)); -- offset MSB 1331
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14632 => state := s14633; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14633 => 			--4
	if (fixed2floatrdy = '1') then state := s14634;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14633; end if;
when s14634 => state := s14635; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14635 => 			--6
	if (mulfprdy = '1') then state := s14636;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14635; end if;
when s14636 => state := s14637; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14637 => 			--8
	if (mulfprdy = '1') then state := s14638;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14637; end if;
when s14638 => state := s14639; 	--9
	mulfpsclr <= '0';
when s14639 => state := s14640; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14640 => 			--11
	if (mulfprdy = '1') then state := s14641;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14640; end if;
when s14641 => state := s14642; 	--12
	mulfpsclr <= '0';
when s14642 => state := s14643; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14643 => 			--14
	if (addfprdy = '1') then state := s14644;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14643; end if;
when s14644 => state := s14645; 	--15
	addfpsclr <= '0';
when s14645 => state := s14646; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14646 => 			--17
	if (addfprdy = '1') then state := s14647;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14646; end if;
when s14647 => state := s14648; 	--18
	addfpsclr <= '0';
when s14648 => state := s14649; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14649 => 			--20
	if (addfprdy = '1') then state := s14650;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14649; end if;
when s14650 => state := s14651; 	--21
	addfpsclr <= '0';
when s14651 => state := s14652; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (721, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14652 => state := s14653; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1380, 12)); -- offset LSB 1332
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s14653 => state := s14654;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1381, 12)); -- offset MSB 1333
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14654 => state := s14655; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14655 => 			--4
	if (fixed2floatrdy = '1') then state := s14656;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14655; end if;
when s14656 => state := s14657; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14657 => 			--6
	if (mulfprdy = '1') then state := s14658;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14657; end if;
when s14658 => state := s14659; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14659 => 			--8
	if (mulfprdy = '1') then state := s14660;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14659; end if;
when s14660 => state := s14661; 	--9
	mulfpsclr <= '0';
when s14661 => state := s14662; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14662 => 			--11
	if (mulfprdy = '1') then state := s14663;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14662; end if;
when s14663 => state := s14664; 	--12
	mulfpsclr <= '0';
when s14664 => state := s14665; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14665 => 			--14
	if (addfprdy = '1') then state := s14666;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14665; end if;
when s14666 => state := s14667; 	--15
	addfpsclr <= '0';
when s14667 => state := s14668; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14668 => 			--17
	if (addfprdy = '1') then state := s14669;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14668; end if;
when s14669 => state := s14670; 	--18
	addfpsclr <= '0';
when s14670 => state := s14671; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14671 => 			--20
	if (addfprdy = '1') then state := s14672;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14671; end if;
when s14672 => state := s14673; 	--21
	addfpsclr <= '0';
when s14673 => state := s14674; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (722, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14674 => state := s14675; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1382, 12)); -- offset LSB 1334
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s14675 => state := s14676;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1383, 12)); -- offset MSB 1335
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14676 => state := s14677; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14677 => 			--4
	if (fixed2floatrdy = '1') then state := s14678;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14677; end if;
when s14678 => state := s14679; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14679 => 			--6
	if (mulfprdy = '1') then state := s14680;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14679; end if;
when s14680 => state := s14681; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14681 => 			--8
	if (mulfprdy = '1') then state := s14682;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14681; end if;
when s14682 => state := s14683; 	--9
	mulfpsclr <= '0';
when s14683 => state := s14684; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14684 => 			--11
	if (mulfprdy = '1') then state := s14685;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14684; end if;
when s14685 => state := s14686; 	--12
	mulfpsclr <= '0';
when s14686 => state := s14687; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14687 => 			--14
	if (addfprdy = '1') then state := s14688;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14687; end if;
when s14688 => state := s14689; 	--15
	addfpsclr <= '0';
when s14689 => state := s14690; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14690 => 			--17
	if (addfprdy = '1') then state := s14691;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14690; end if;
when s14691 => state := s14692; 	--18
	addfpsclr <= '0';
when s14692 => state := s14693; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14693 => 			--20
	if (addfprdy = '1') then state := s14694;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14693; end if;
when s14694 => state := s14695; 	--21
	addfpsclr <= '0';
when s14695 => state := s14696; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (723, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14696 => state := s14697; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1384, 12)); -- offset LSB 1336
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s14697 => state := s14698;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1385, 12)); -- offset MSB 1337
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14698 => state := s14699; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14699 => 			--4
	if (fixed2floatrdy = '1') then state := s14700;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14699; end if;
when s14700 => state := s14701; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14701 => 			--6
	if (mulfprdy = '1') then state := s14702;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14701; end if;
when s14702 => state := s14703; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14703 => 			--8
	if (mulfprdy = '1') then state := s14704;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14703; end if;
when s14704 => state := s14705; 	--9
	mulfpsclr <= '0';
when s14705 => state := s14706; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14706 => 			--11
	if (mulfprdy = '1') then state := s14707;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14706; end if;
when s14707 => state := s14708; 	--12
	mulfpsclr <= '0';
when s14708 => state := s14709; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14709 => 			--14
	if (addfprdy = '1') then state := s14710;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14709; end if;
when s14710 => state := s14711; 	--15
	addfpsclr <= '0';
when s14711 => state := s14712; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14712 => 			--17
	if (addfprdy = '1') then state := s14713;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14712; end if;
when s14713 => state := s14714; 	--18
	addfpsclr <= '0';
when s14714 => state := s14715; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14715 => 			--20
	if (addfprdy = '1') then state := s14716;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14715; end if;
when s14716 => state := s14717; 	--21
	addfpsclr <= '0';
when s14717 => state := s14718; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (724, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14718 => state := s14719; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1386, 12)); -- offset LSB 1338
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s14719 => state := s14720;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1387, 12)); -- offset MSB 1339
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14720 => state := s14721; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14721 => 			--4
	if (fixed2floatrdy = '1') then state := s14722;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14721; end if;
when s14722 => state := s14723; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14723 => 			--6
	if (mulfprdy = '1') then state := s14724;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14723; end if;
when s14724 => state := s14725; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14725 => 			--8
	if (mulfprdy = '1') then state := s14726;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14725; end if;
when s14726 => state := s14727; 	--9
	mulfpsclr <= '0';
when s14727 => state := s14728; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14728 => 			--11
	if (mulfprdy = '1') then state := s14729;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14728; end if;
when s14729 => state := s14730; 	--12
	mulfpsclr <= '0';
when s14730 => state := s14731; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14731 => 			--14
	if (addfprdy = '1') then state := s14732;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14731; end if;
when s14732 => state := s14733; 	--15
	addfpsclr <= '0';
when s14733 => state := s14734; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14734 => 			--17
	if (addfprdy = '1') then state := s14735;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14734; end if;
when s14735 => state := s14736; 	--18
	addfpsclr <= '0';
when s14736 => state := s14737; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14737 => 			--20
	if (addfprdy = '1') then state := s14738;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14737; end if;
when s14738 => state := s14739; 	--21
	addfpsclr <= '0';
when s14739 => state := s14740; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (725, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14740 => state := s14741; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1388, 12)); -- offset LSB 1340
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s14741 => state := s14742;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1389, 12)); -- offset MSB 1341
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14742 => state := s14743; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14743 => 			--4
	if (fixed2floatrdy = '1') then state := s14744;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14743; end if;
when s14744 => state := s14745; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14745 => 			--6
	if (mulfprdy = '1') then state := s14746;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14745; end if;
when s14746 => state := s14747; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14747 => 			--8
	if (mulfprdy = '1') then state := s14748;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14747; end if;
when s14748 => state := s14749; 	--9
	mulfpsclr <= '0';
when s14749 => state := s14750; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14750 => 			--11
	if (mulfprdy = '1') then state := s14751;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14750; end if;
when s14751 => state := s14752; 	--12
	mulfpsclr <= '0';
when s14752 => state := s14753; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14753 => 			--14
	if (addfprdy = '1') then state := s14754;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14753; end if;
when s14754 => state := s14755; 	--15
	addfpsclr <= '0';
when s14755 => state := s14756; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14756 => 			--17
	if (addfprdy = '1') then state := s14757;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14756; end if;
when s14757 => state := s14758; 	--18
	addfpsclr <= '0';
when s14758 => state := s14759; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14759 => 			--20
	if (addfprdy = '1') then state := s14760;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14759; end if;
when s14760 => state := s14761; 	--21
	addfpsclr <= '0';
when s14761 => state := s14762; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (726, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14762 => state := s14763; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1390, 12)); -- offset LSB 1342
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s14763 => state := s14764;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1391, 12)); -- offset MSB 1343
	addra <= std_logic_vector (to_unsigned (20, 10)); -- OCCrowI 20
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14764 => state := s14765; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14765 => 			--4
	if (fixed2floatrdy = '1') then state := s14766;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14765; end if;
when s14766 => state := s14767; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14767 => 			--6
	if (mulfprdy = '1') then state := s14768;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14767; end if;
when s14768 => state := s14769; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14769 => 			--8
	if (mulfprdy = '1') then state := s14770;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14769; end if;
when s14770 => state := s14771; 	--9
	mulfpsclr <= '0';
when s14771 => state := s14772; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14772 => 			--11
	if (mulfprdy = '1') then state := s14773;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14772; end if;
when s14773 => state := s14774; 	--12
	mulfpsclr <= '0';
when s14774 => state := s14775; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14775 => 			--14
	if (addfprdy = '1') then state := s14776;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14775; end if;
when s14776 => state := s14777; 	--15
	addfpsclr <= '0';
when s14777 => state := s14778; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14778 => 			--17
	if (addfprdy = '1') then state := s14779;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14778; end if;
when s14779 => state := s14780; 	--18
	addfpsclr <= '0';
when s14780 => state := s14781; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14781 => 			--20
	if (addfprdy = '1') then state := s14782;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14781; end if;
when s14782 => state := s14783; 	--21
	addfpsclr <= '0';
when s14783 => state := s14784; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (727, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14784 => state := s14785; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1392, 12)); -- offset LSB 1344
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s14785 => state := s14786;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1393, 12)); -- offset MSB 1345
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14786 => state := s14787; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14787 => 			--4
	if (fixed2floatrdy = '1') then state := s14788;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14787; end if;
when s14788 => state := s14789; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14789 => 			--6
	if (mulfprdy = '1') then state := s14790;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14789; end if;
when s14790 => state := s14791; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14791 => 			--8
	if (mulfprdy = '1') then state := s14792;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14791; end if;
when s14792 => state := s14793; 	--9
	mulfpsclr <= '0';
when s14793 => state := s14794; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14794 => 			--11
	if (mulfprdy = '1') then state := s14795;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14794; end if;
when s14795 => state := s14796; 	--12
	mulfpsclr <= '0';
when s14796 => state := s14797; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14797 => 			--14
	if (addfprdy = '1') then state := s14798;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14797; end if;
when s14798 => state := s14799; 	--15
	addfpsclr <= '0';
when s14799 => state := s14800; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14800 => 			--17
	if (addfprdy = '1') then state := s14801;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14800; end if;
when s14801 => state := s14802; 	--18
	addfpsclr <= '0';
when s14802 => state := s14803; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14803 => 			--20
	if (addfprdy = '1') then state := s14804;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14803; end if;
when s14804 => state := s14805; 	--21
	addfpsclr <= '0';
when s14805 => state := s14806; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (728, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14806 => state := s14807; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1394, 12)); -- offset LSB 1346
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s14807 => state := s14808;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1395, 12)); -- offset MSB 1347
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14808 => state := s14809; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14809 => 			--4
	if (fixed2floatrdy = '1') then state := s14810;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14809; end if;
when s14810 => state := s14811; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14811 => 			--6
	if (mulfprdy = '1') then state := s14812;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14811; end if;
when s14812 => state := s14813; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14813 => 			--8
	if (mulfprdy = '1') then state := s14814;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14813; end if;
when s14814 => state := s14815; 	--9
	mulfpsclr <= '0';
when s14815 => state := s14816; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14816 => 			--11
	if (mulfprdy = '1') then state := s14817;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14816; end if;
when s14817 => state := s14818; 	--12
	mulfpsclr <= '0';
when s14818 => state := s14819; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14819 => 			--14
	if (addfprdy = '1') then state := s14820;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14819; end if;
when s14820 => state := s14821; 	--15
	addfpsclr <= '0';
when s14821 => state := s14822; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14822 => 			--17
	if (addfprdy = '1') then state := s14823;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14822; end if;
when s14823 => state := s14824; 	--18
	addfpsclr <= '0';
when s14824 => state := s14825; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14825 => 			--20
	if (addfprdy = '1') then state := s14826;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14825; end if;
when s14826 => state := s14827; 	--21
	addfpsclr <= '0';
when s14827 => state := s14828; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (729, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14828 => state := s14829; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1396, 12)); -- offset LSB 1348
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s14829 => state := s14830;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1397, 12)); -- offset MSB 1349
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14830 => state := s14831; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14831 => 			--4
	if (fixed2floatrdy = '1') then state := s14832;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14831; end if;
when s14832 => state := s14833; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14833 => 			--6
	if (mulfprdy = '1') then state := s14834;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14833; end if;
when s14834 => state := s14835; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14835 => 			--8
	if (mulfprdy = '1') then state := s14836;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14835; end if;
when s14836 => state := s14837; 	--9
	mulfpsclr <= '0';
when s14837 => state := s14838; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14838 => 			--11
	if (mulfprdy = '1') then state := s14839;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14838; end if;
when s14839 => state := s14840; 	--12
	mulfpsclr <= '0';
when s14840 => state := s14841; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14841 => 			--14
	if (addfprdy = '1') then state := s14842;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14841; end if;
when s14842 => state := s14843; 	--15
	addfpsclr <= '0';
when s14843 => state := s14844; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14844 => 			--17
	if (addfprdy = '1') then state := s14845;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14844; end if;
when s14845 => state := s14846; 	--18
	addfpsclr <= '0';
when s14846 => state := s14847; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14847 => 			--20
	if (addfprdy = '1') then state := s14848;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14847; end if;
when s14848 => state := s14849; 	--21
	addfpsclr <= '0';
when s14849 => state := s14850; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (730, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14850 => state := s14851; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1398, 12)); -- offset LSB 1350
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s14851 => state := s14852;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1399, 12)); -- offset MSB 1351
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14852 => state := s14853; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14853 => 			--4
	if (fixed2floatrdy = '1') then state := s14854;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14853; end if;
when s14854 => state := s14855; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14855 => 			--6
	if (mulfprdy = '1') then state := s14856;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14855; end if;
when s14856 => state := s14857; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14857 => 			--8
	if (mulfprdy = '1') then state := s14858;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14857; end if;
when s14858 => state := s14859; 	--9
	mulfpsclr <= '0';
when s14859 => state := s14860; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14860 => 			--11
	if (mulfprdy = '1') then state := s14861;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14860; end if;
when s14861 => state := s14862; 	--12
	mulfpsclr <= '0';
when s14862 => state := s14863; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14863 => 			--14
	if (addfprdy = '1') then state := s14864;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14863; end if;
when s14864 => state := s14865; 	--15
	addfpsclr <= '0';
when s14865 => state := s14866; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14866 => 			--17
	if (addfprdy = '1') then state := s14867;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14866; end if;
when s14867 => state := s14868; 	--18
	addfpsclr <= '0';
when s14868 => state := s14869; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14869 => 			--20
	if (addfprdy = '1') then state := s14870;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14869; end if;
when s14870 => state := s14871; 	--21
	addfpsclr <= '0';
when s14871 => state := s14872; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (731, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14872 => state := s14873; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1400, 12)); -- offset LSB 1352
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s14873 => state := s14874;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1401, 12)); -- offset MSB 1353
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14874 => state := s14875; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14875 => 			--4
	if (fixed2floatrdy = '1') then state := s14876;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14875; end if;
when s14876 => state := s14877; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14877 => 			--6
	if (mulfprdy = '1') then state := s14878;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14877; end if;
when s14878 => state := s14879; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14879 => 			--8
	if (mulfprdy = '1') then state := s14880;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14879; end if;
when s14880 => state := s14881; 	--9
	mulfpsclr <= '0';
when s14881 => state := s14882; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14882 => 			--11
	if (mulfprdy = '1') then state := s14883;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14882; end if;
when s14883 => state := s14884; 	--12
	mulfpsclr <= '0';
when s14884 => state := s14885; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14885 => 			--14
	if (addfprdy = '1') then state := s14886;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14885; end if;
when s14886 => state := s14887; 	--15
	addfpsclr <= '0';
when s14887 => state := s14888; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14888 => 			--17
	if (addfprdy = '1') then state := s14889;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14888; end if;
when s14889 => state := s14890; 	--18
	addfpsclr <= '0';
when s14890 => state := s14891; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14891 => 			--20
	if (addfprdy = '1') then state := s14892;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14891; end if;
when s14892 => state := s14893; 	--21
	addfpsclr <= '0';
when s14893 => state := s14894; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (732, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14894 => state := s14895; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1402, 12)); -- offset LSB 1354
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s14895 => state := s14896;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1403, 12)); -- offset MSB 1355
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14896 => state := s14897; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14897 => 			--4
	if (fixed2floatrdy = '1') then state := s14898;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14897; end if;
when s14898 => state := s14899; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14899 => 			--6
	if (mulfprdy = '1') then state := s14900;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14899; end if;
when s14900 => state := s14901; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14901 => 			--8
	if (mulfprdy = '1') then state := s14902;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14901; end if;
when s14902 => state := s14903; 	--9
	mulfpsclr <= '0';
when s14903 => state := s14904; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14904 => 			--11
	if (mulfprdy = '1') then state := s14905;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14904; end if;
when s14905 => state := s14906; 	--12
	mulfpsclr <= '0';
when s14906 => state := s14907; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14907 => 			--14
	if (addfprdy = '1') then state := s14908;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14907; end if;
when s14908 => state := s14909; 	--15
	addfpsclr <= '0';
when s14909 => state := s14910; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14910 => 			--17
	if (addfprdy = '1') then state := s14911;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14910; end if;
when s14911 => state := s14912; 	--18
	addfpsclr <= '0';
when s14912 => state := s14913; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14913 => 			--20
	if (addfprdy = '1') then state := s14914;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14913; end if;
when s14914 => state := s14915; 	--21
	addfpsclr <= '0';
when s14915 => state := s14916; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (733, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14916 => state := s14917; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1404, 12)); -- offset LSB 1356
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s14917 => state := s14918;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1405, 12)); -- offset MSB 1357
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14918 => state := s14919; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14919 => 			--4
	if (fixed2floatrdy = '1') then state := s14920;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14919; end if;
when s14920 => state := s14921; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14921 => 			--6
	if (mulfprdy = '1') then state := s14922;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14921; end if;
when s14922 => state := s14923; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14923 => 			--8
	if (mulfprdy = '1') then state := s14924;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14923; end if;
when s14924 => state := s14925; 	--9
	mulfpsclr <= '0';
when s14925 => state := s14926; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14926 => 			--11
	if (mulfprdy = '1') then state := s14927;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14926; end if;
when s14927 => state := s14928; 	--12
	mulfpsclr <= '0';
when s14928 => state := s14929; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14929 => 			--14
	if (addfprdy = '1') then state := s14930;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14929; end if;
when s14930 => state := s14931; 	--15
	addfpsclr <= '0';
when s14931 => state := s14932; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14932 => 			--17
	if (addfprdy = '1') then state := s14933;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14932; end if;
when s14933 => state := s14934; 	--18
	addfpsclr <= '0';
when s14934 => state := s14935; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14935 => 			--20
	if (addfprdy = '1') then state := s14936;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14935; end if;
when s14936 => state := s14937; 	--21
	addfpsclr <= '0';
when s14937 => state := s14938; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (734, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14938 => state := s14939; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1406, 12)); -- offset LSB 1358
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s14939 => state := s14940;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1407, 12)); -- offset MSB 1359
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14940 => state := s14941; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14941 => 			--4
	if (fixed2floatrdy = '1') then state := s14942;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14941; end if;
when s14942 => state := s14943; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14943 => 			--6
	if (mulfprdy = '1') then state := s14944;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14943; end if;
when s14944 => state := s14945; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14945 => 			--8
	if (mulfprdy = '1') then state := s14946;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14945; end if;
when s14946 => state := s14947; 	--9
	mulfpsclr <= '0';
when s14947 => state := s14948; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14948 => 			--11
	if (mulfprdy = '1') then state := s14949;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14948; end if;
when s14949 => state := s14950; 	--12
	mulfpsclr <= '0';
when s14950 => state := s14951; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14951 => 			--14
	if (addfprdy = '1') then state := s14952;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14951; end if;
when s14952 => state := s14953; 	--15
	addfpsclr <= '0';
when s14953 => state := s14954; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14954 => 			--17
	if (addfprdy = '1') then state := s14955;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14954; end if;
when s14955 => state := s14956; 	--18
	addfpsclr <= '0';
when s14956 => state := s14957; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14957 => 			--20
	if (addfprdy = '1') then state := s14958;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14957; end if;
when s14958 => state := s14959; 	--21
	addfpsclr <= '0';
when s14959 => state := s14960; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (735, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14960 => state := s14961; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1408, 12)); -- offset LSB 1360
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s14961 => state := s14962;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1409, 12)); -- offset MSB 1361
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14962 => state := s14963; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14963 => 			--4
	if (fixed2floatrdy = '1') then state := s14964;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14963; end if;
when s14964 => state := s14965; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14965 => 			--6
	if (mulfprdy = '1') then state := s14966;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14965; end if;
when s14966 => state := s14967; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14967 => 			--8
	if (mulfprdy = '1') then state := s14968;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14967; end if;
when s14968 => state := s14969; 	--9
	mulfpsclr <= '0';
when s14969 => state := s14970; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14970 => 			--11
	if (mulfprdy = '1') then state := s14971;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14970; end if;
when s14971 => state := s14972; 	--12
	mulfpsclr <= '0';
when s14972 => state := s14973; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14973 => 			--14
	if (addfprdy = '1') then state := s14974;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14973; end if;
when s14974 => state := s14975; 	--15
	addfpsclr <= '0';
when s14975 => state := s14976; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14976 => 			--17
	if (addfprdy = '1') then state := s14977;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14976; end if;
when s14977 => state := s14978; 	--18
	addfpsclr <= '0';
when s14978 => state := s14979; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s14979 => 			--20
	if (addfprdy = '1') then state := s14980;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14979; end if;
when s14980 => state := s14981; 	--21
	addfpsclr <= '0';
when s14981 => state := s14982; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (736, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s14982 => state := s14983; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1410, 12)); -- offset LSB 1362
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s14983 => state := s14984;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1411, 12)); -- offset MSB 1363
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s14984 => state := s14985; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s14985 => 			--4
	if (fixed2floatrdy = '1') then state := s14986;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s14985; end if;
when s14986 => state := s14987; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s14987 => 			--6
	if (mulfprdy = '1') then state := s14988;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14987; end if;
when s14988 => state := s14989; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s14989 => 			--8
	if (mulfprdy = '1') then state := s14990;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14989; end if;
when s14990 => state := s14991; 	--9
	mulfpsclr <= '0';
when s14991 => state := s14992; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s14992 => 			--11
	if (mulfprdy = '1') then state := s14993;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s14992; end if;
when s14993 => state := s14994; 	--12
	mulfpsclr <= '0';
when s14994 => state := s14995; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s14995 => 			--14
	if (addfprdy = '1') then state := s14996;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14995; end if;
when s14996 => state := s14997; 	--15
	addfpsclr <= '0';
when s14997 => state := s14998; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s14998 => 			--17
	if (addfprdy = '1') then state := s14999;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s14998; end if;
when s14999 => state := s15000; 	--18
	addfpsclr <= '0';
when s15000 => state := s15001; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15001 => 			--20
	if (addfprdy = '1') then state := s15002;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15001; end if;
when s15002 => state := s15003; 	--21
	addfpsclr <= '0';
when s15003 => state := s15004; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (737, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15004 => state := s15005; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1412, 12)); -- offset LSB 1364
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s15005 => state := s15006;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1413, 12)); -- offset MSB 1365
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15006 => state := s15007; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15007 => 			--4
	if (fixed2floatrdy = '1') then state := s15008;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15007; end if;
when s15008 => state := s15009; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15009 => 			--6
	if (mulfprdy = '1') then state := s15010;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15009; end if;
when s15010 => state := s15011; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15011 => 			--8
	if (mulfprdy = '1') then state := s15012;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15011; end if;
when s15012 => state := s15013; 	--9
	mulfpsclr <= '0';
when s15013 => state := s15014; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15014 => 			--11
	if (mulfprdy = '1') then state := s15015;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15014; end if;
when s15015 => state := s15016; 	--12
	mulfpsclr <= '0';
when s15016 => state := s15017; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15017 => 			--14
	if (addfprdy = '1') then state := s15018;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15017; end if;
when s15018 => state := s15019; 	--15
	addfpsclr <= '0';
when s15019 => state := s15020; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15020 => 			--17
	if (addfprdy = '1') then state := s15021;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15020; end if;
when s15021 => state := s15022; 	--18
	addfpsclr <= '0';
when s15022 => state := s15023; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15023 => 			--20
	if (addfprdy = '1') then state := s15024;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15023; end if;
when s15024 => state := s15025; 	--21
	addfpsclr <= '0';
when s15025 => state := s15026; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (738, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15026 => state := s15027; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1414, 12)); -- offset LSB 1366
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s15027 => state := s15028;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1415, 12)); -- offset MSB 1367
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15028 => state := s15029; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15029 => 			--4
	if (fixed2floatrdy = '1') then state := s15030;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15029; end if;
when s15030 => state := s15031; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15031 => 			--6
	if (mulfprdy = '1') then state := s15032;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15031; end if;
when s15032 => state := s15033; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15033 => 			--8
	if (mulfprdy = '1') then state := s15034;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15033; end if;
when s15034 => state := s15035; 	--9
	mulfpsclr <= '0';
when s15035 => state := s15036; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15036 => 			--11
	if (mulfprdy = '1') then state := s15037;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15036; end if;
when s15037 => state := s15038; 	--12
	mulfpsclr <= '0';
when s15038 => state := s15039; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15039 => 			--14
	if (addfprdy = '1') then state := s15040;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15039; end if;
when s15040 => state := s15041; 	--15
	addfpsclr <= '0';
when s15041 => state := s15042; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15042 => 			--17
	if (addfprdy = '1') then state := s15043;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15042; end if;
when s15043 => state := s15044; 	--18
	addfpsclr <= '0';
when s15044 => state := s15045; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15045 => 			--20
	if (addfprdy = '1') then state := s15046;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15045; end if;
when s15046 => state := s15047; 	--21
	addfpsclr <= '0';
when s15047 => state := s15048; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (739, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15048 => state := s15049; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1416, 12)); -- offset LSB 1368
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s15049 => state := s15050;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1417, 12)); -- offset MSB 1369
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15050 => state := s15051; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15051 => 			--4
	if (fixed2floatrdy = '1') then state := s15052;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15051; end if;
when s15052 => state := s15053; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15053 => 			--6
	if (mulfprdy = '1') then state := s15054;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15053; end if;
when s15054 => state := s15055; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15055 => 			--8
	if (mulfprdy = '1') then state := s15056;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15055; end if;
when s15056 => state := s15057; 	--9
	mulfpsclr <= '0';
when s15057 => state := s15058; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15058 => 			--11
	if (mulfprdy = '1') then state := s15059;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15058; end if;
when s15059 => state := s15060; 	--12
	mulfpsclr <= '0';
when s15060 => state := s15061; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15061 => 			--14
	if (addfprdy = '1') then state := s15062;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15061; end if;
when s15062 => state := s15063; 	--15
	addfpsclr <= '0';
when s15063 => state := s15064; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15064 => 			--17
	if (addfprdy = '1') then state := s15065;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15064; end if;
when s15065 => state := s15066; 	--18
	addfpsclr <= '0';
when s15066 => state := s15067; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15067 => 			--20
	if (addfprdy = '1') then state := s15068;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15067; end if;
when s15068 => state := s15069; 	--21
	addfpsclr <= '0';
when s15069 => state := s15070; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (740, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15070 => state := s15071; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1418, 12)); -- offset LSB 1370
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s15071 => state := s15072;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1419, 12)); -- offset MSB 1371
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15072 => state := s15073; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15073 => 			--4
	if (fixed2floatrdy = '1') then state := s15074;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15073; end if;
when s15074 => state := s15075; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15075 => 			--6
	if (mulfprdy = '1') then state := s15076;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15075; end if;
when s15076 => state := s15077; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15077 => 			--8
	if (mulfprdy = '1') then state := s15078;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15077; end if;
when s15078 => state := s15079; 	--9
	mulfpsclr <= '0';
when s15079 => state := s15080; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15080 => 			--11
	if (mulfprdy = '1') then state := s15081;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15080; end if;
when s15081 => state := s15082; 	--12
	mulfpsclr <= '0';
when s15082 => state := s15083; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15083 => 			--14
	if (addfprdy = '1') then state := s15084;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15083; end if;
when s15084 => state := s15085; 	--15
	addfpsclr <= '0';
when s15085 => state := s15086; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15086 => 			--17
	if (addfprdy = '1') then state := s15087;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15086; end if;
when s15087 => state := s15088; 	--18
	addfpsclr <= '0';
when s15088 => state := s15089; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15089 => 			--20
	if (addfprdy = '1') then state := s15090;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15089; end if;
when s15090 => state := s15091; 	--21
	addfpsclr <= '0';
when s15091 => state := s15092; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (741, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15092 => state := s15093; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1420, 12)); -- offset LSB 1372
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s15093 => state := s15094;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1421, 12)); -- offset MSB 1373
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15094 => state := s15095; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15095 => 			--4
	if (fixed2floatrdy = '1') then state := s15096;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15095; end if;
when s15096 => state := s15097; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15097 => 			--6
	if (mulfprdy = '1') then state := s15098;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15097; end if;
when s15098 => state := s15099; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15099 => 			--8
	if (mulfprdy = '1') then state := s15100;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15099; end if;
when s15100 => state := s15101; 	--9
	mulfpsclr <= '0';
when s15101 => state := s15102; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15102 => 			--11
	if (mulfprdy = '1') then state := s15103;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15102; end if;
when s15103 => state := s15104; 	--12
	mulfpsclr <= '0';
when s15104 => state := s15105; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15105 => 			--14
	if (addfprdy = '1') then state := s15106;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15105; end if;
when s15106 => state := s15107; 	--15
	addfpsclr <= '0';
when s15107 => state := s15108; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15108 => 			--17
	if (addfprdy = '1') then state := s15109;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15108; end if;
when s15109 => state := s15110; 	--18
	addfpsclr <= '0';
when s15110 => state := s15111; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15111 => 			--20
	if (addfprdy = '1') then state := s15112;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15111; end if;
when s15112 => state := s15113; 	--21
	addfpsclr <= '0';
when s15113 => state := s15114; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (742, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15114 => state := s15115; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1422, 12)); -- offset LSB 1374
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s15115 => state := s15116;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1423, 12)); -- offset MSB 1375
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15116 => state := s15117; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15117 => 			--4
	if (fixed2floatrdy = '1') then state := s15118;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15117; end if;
when s15118 => state := s15119; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15119 => 			--6
	if (mulfprdy = '1') then state := s15120;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15119; end if;
when s15120 => state := s15121; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15121 => 			--8
	if (mulfprdy = '1') then state := s15122;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15121; end if;
when s15122 => state := s15123; 	--9
	mulfpsclr <= '0';
when s15123 => state := s15124; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15124 => 			--11
	if (mulfprdy = '1') then state := s15125;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15124; end if;
when s15125 => state := s15126; 	--12
	mulfpsclr <= '0';
when s15126 => state := s15127; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15127 => 			--14
	if (addfprdy = '1') then state := s15128;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15127; end if;
when s15128 => state := s15129; 	--15
	addfpsclr <= '0';
when s15129 => state := s15130; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15130 => 			--17
	if (addfprdy = '1') then state := s15131;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15130; end if;
when s15131 => state := s15132; 	--18
	addfpsclr <= '0';
when s15132 => state := s15133; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15133 => 			--20
	if (addfprdy = '1') then state := s15134;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15133; end if;
when s15134 => state := s15135; 	--21
	addfpsclr <= '0';
when s15135 => state := s15136; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (743, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15136 => state := s15137; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1424, 12)); -- offset LSB 1376
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s15137 => state := s15138;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1425, 12)); -- offset MSB 1377
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15138 => state := s15139; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15139 => 			--4
	if (fixed2floatrdy = '1') then state := s15140;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15139; end if;
when s15140 => state := s15141; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15141 => 			--6
	if (mulfprdy = '1') then state := s15142;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15141; end if;
when s15142 => state := s15143; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15143 => 			--8
	if (mulfprdy = '1') then state := s15144;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15143; end if;
when s15144 => state := s15145; 	--9
	mulfpsclr <= '0';
when s15145 => state := s15146; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15146 => 			--11
	if (mulfprdy = '1') then state := s15147;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15146; end if;
when s15147 => state := s15148; 	--12
	mulfpsclr <= '0';
when s15148 => state := s15149; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15149 => 			--14
	if (addfprdy = '1') then state := s15150;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15149; end if;
when s15150 => state := s15151; 	--15
	addfpsclr <= '0';
when s15151 => state := s15152; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15152 => 			--17
	if (addfprdy = '1') then state := s15153;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15152; end if;
when s15153 => state := s15154; 	--18
	addfpsclr <= '0';
when s15154 => state := s15155; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15155 => 			--20
	if (addfprdy = '1') then state := s15156;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15155; end if;
when s15156 => state := s15157; 	--21
	addfpsclr <= '0';
when s15157 => state := s15158; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (744, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15158 => state := s15159; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1426, 12)); -- offset LSB 1378
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s15159 => state := s15160;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1427, 12)); -- offset MSB 1379
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15160 => state := s15161; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15161 => 			--4
	if (fixed2floatrdy = '1') then state := s15162;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15161; end if;
when s15162 => state := s15163; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15163 => 			--6
	if (mulfprdy = '1') then state := s15164;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15163; end if;
when s15164 => state := s15165; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15165 => 			--8
	if (mulfprdy = '1') then state := s15166;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15165; end if;
when s15166 => state := s15167; 	--9
	mulfpsclr <= '0';
when s15167 => state := s15168; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15168 => 			--11
	if (mulfprdy = '1') then state := s15169;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15168; end if;
when s15169 => state := s15170; 	--12
	mulfpsclr <= '0';
when s15170 => state := s15171; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15171 => 			--14
	if (addfprdy = '1') then state := s15172;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15171; end if;
when s15172 => state := s15173; 	--15
	addfpsclr <= '0';
when s15173 => state := s15174; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15174 => 			--17
	if (addfprdy = '1') then state := s15175;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15174; end if;
when s15175 => state := s15176; 	--18
	addfpsclr <= '0';
when s15176 => state := s15177; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15177 => 			--20
	if (addfprdy = '1') then state := s15178;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15177; end if;
when s15178 => state := s15179; 	--21
	addfpsclr <= '0';
when s15179 => state := s15180; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (745, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15180 => state := s15181; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1428, 12)); -- offset LSB 1380
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s15181 => state := s15182;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1429, 12)); -- offset MSB 1381
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15182 => state := s15183; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15183 => 			--4
	if (fixed2floatrdy = '1') then state := s15184;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15183; end if;
when s15184 => state := s15185; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15185 => 			--6
	if (mulfprdy = '1') then state := s15186;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15185; end if;
when s15186 => state := s15187; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15187 => 			--8
	if (mulfprdy = '1') then state := s15188;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15187; end if;
when s15188 => state := s15189; 	--9
	mulfpsclr <= '0';
when s15189 => state := s15190; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15190 => 			--11
	if (mulfprdy = '1') then state := s15191;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15190; end if;
when s15191 => state := s15192; 	--12
	mulfpsclr <= '0';
when s15192 => state := s15193; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15193 => 			--14
	if (addfprdy = '1') then state := s15194;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15193; end if;
when s15194 => state := s15195; 	--15
	addfpsclr <= '0';
when s15195 => state := s15196; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15196 => 			--17
	if (addfprdy = '1') then state := s15197;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15196; end if;
when s15197 => state := s15198; 	--18
	addfpsclr <= '0';
when s15198 => state := s15199; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15199 => 			--20
	if (addfprdy = '1') then state := s15200;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15199; end if;
when s15200 => state := s15201; 	--21
	addfpsclr <= '0';
when s15201 => state := s15202; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (746, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15202 => state := s15203; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1430, 12)); -- offset LSB 1382
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s15203 => state := s15204;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1431, 12)); -- offset MSB 1383
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15204 => state := s15205; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15205 => 			--4
	if (fixed2floatrdy = '1') then state := s15206;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15205; end if;
when s15206 => state := s15207; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15207 => 			--6
	if (mulfprdy = '1') then state := s15208;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15207; end if;
when s15208 => state := s15209; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15209 => 			--8
	if (mulfprdy = '1') then state := s15210;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15209; end if;
when s15210 => state := s15211; 	--9
	mulfpsclr <= '0';
when s15211 => state := s15212; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15212 => 			--11
	if (mulfprdy = '1') then state := s15213;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15212; end if;
when s15213 => state := s15214; 	--12
	mulfpsclr <= '0';
when s15214 => state := s15215; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15215 => 			--14
	if (addfprdy = '1') then state := s15216;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15215; end if;
when s15216 => state := s15217; 	--15
	addfpsclr <= '0';
when s15217 => state := s15218; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15218 => 			--17
	if (addfprdy = '1') then state := s15219;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15218; end if;
when s15219 => state := s15220; 	--18
	addfpsclr <= '0';
when s15220 => state := s15221; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15221 => 			--20
	if (addfprdy = '1') then state := s15222;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15221; end if;
when s15222 => state := s15223; 	--21
	addfpsclr <= '0';
when s15223 => state := s15224; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (747, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15224 => state := s15225; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1432, 12)); -- offset LSB 1384
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s15225 => state := s15226;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1433, 12)); -- offset MSB 1385
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15226 => state := s15227; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15227 => 			--4
	if (fixed2floatrdy = '1') then state := s15228;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15227; end if;
when s15228 => state := s15229; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15229 => 			--6
	if (mulfprdy = '1') then state := s15230;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15229; end if;
when s15230 => state := s15231; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15231 => 			--8
	if (mulfprdy = '1') then state := s15232;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15231; end if;
when s15232 => state := s15233; 	--9
	mulfpsclr <= '0';
when s15233 => state := s15234; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15234 => 			--11
	if (mulfprdy = '1') then state := s15235;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15234; end if;
when s15235 => state := s15236; 	--12
	mulfpsclr <= '0';
when s15236 => state := s15237; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15237 => 			--14
	if (addfprdy = '1') then state := s15238;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15237; end if;
when s15238 => state := s15239; 	--15
	addfpsclr <= '0';
when s15239 => state := s15240; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15240 => 			--17
	if (addfprdy = '1') then state := s15241;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15240; end if;
when s15241 => state := s15242; 	--18
	addfpsclr <= '0';
when s15242 => state := s15243; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15243 => 			--20
	if (addfprdy = '1') then state := s15244;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15243; end if;
when s15244 => state := s15245; 	--21
	addfpsclr <= '0';
when s15245 => state := s15246; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (748, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15246 => state := s15247; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1434, 12)); -- offset LSB 1386
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s15247 => state := s15248;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1435, 12)); -- offset MSB 1387
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15248 => state := s15249; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15249 => 			--4
	if (fixed2floatrdy = '1') then state := s15250;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15249; end if;
when s15250 => state := s15251; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15251 => 			--6
	if (mulfprdy = '1') then state := s15252;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15251; end if;
when s15252 => state := s15253; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15253 => 			--8
	if (mulfprdy = '1') then state := s15254;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15253; end if;
when s15254 => state := s15255; 	--9
	mulfpsclr <= '0';
when s15255 => state := s15256; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15256 => 			--11
	if (mulfprdy = '1') then state := s15257;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15256; end if;
when s15257 => state := s15258; 	--12
	mulfpsclr <= '0';
when s15258 => state := s15259; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15259 => 			--14
	if (addfprdy = '1') then state := s15260;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15259; end if;
when s15260 => state := s15261; 	--15
	addfpsclr <= '0';
when s15261 => state := s15262; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15262 => 			--17
	if (addfprdy = '1') then state := s15263;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15262; end if;
when s15263 => state := s15264; 	--18
	addfpsclr <= '0';
when s15264 => state := s15265; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15265 => 			--20
	if (addfprdy = '1') then state := s15266;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15265; end if;
when s15266 => state := s15267; 	--21
	addfpsclr <= '0';
when s15267 => state := s15268; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (749, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15268 => state := s15269; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1436, 12)); -- offset LSB 1388
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s15269 => state := s15270;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1437, 12)); -- offset MSB 1389
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15270 => state := s15271; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15271 => 			--4
	if (fixed2floatrdy = '1') then state := s15272;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15271; end if;
when s15272 => state := s15273; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15273 => 			--6
	if (mulfprdy = '1') then state := s15274;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15273; end if;
when s15274 => state := s15275; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15275 => 			--8
	if (mulfprdy = '1') then state := s15276;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15275; end if;
when s15276 => state := s15277; 	--9
	mulfpsclr <= '0';
when s15277 => state := s15278; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15278 => 			--11
	if (mulfprdy = '1') then state := s15279;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15278; end if;
when s15279 => state := s15280; 	--12
	mulfpsclr <= '0';
when s15280 => state := s15281; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15281 => 			--14
	if (addfprdy = '1') then state := s15282;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15281; end if;
when s15282 => state := s15283; 	--15
	addfpsclr <= '0';
when s15283 => state := s15284; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15284 => 			--17
	if (addfprdy = '1') then state := s15285;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15284; end if;
when s15285 => state := s15286; 	--18
	addfpsclr <= '0';
when s15286 => state := s15287; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15287 => 			--20
	if (addfprdy = '1') then state := s15288;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15287; end if;
when s15288 => state := s15289; 	--21
	addfpsclr <= '0';
when s15289 => state := s15290; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (750, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15290 => state := s15291; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1438, 12)); -- offset LSB 1390
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s15291 => state := s15292;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1439, 12)); -- offset MSB 1391
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15292 => state := s15293; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15293 => 			--4
	if (fixed2floatrdy = '1') then state := s15294;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15293; end if;
when s15294 => state := s15295; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15295 => 			--6
	if (mulfprdy = '1') then state := s15296;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15295; end if;
when s15296 => state := s15297; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15297 => 			--8
	if (mulfprdy = '1') then state := s15298;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15297; end if;
when s15298 => state := s15299; 	--9
	mulfpsclr <= '0';
when s15299 => state := s15300; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15300 => 			--11
	if (mulfprdy = '1') then state := s15301;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15300; end if;
when s15301 => state := s15302; 	--12
	mulfpsclr <= '0';
when s15302 => state := s15303; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15303 => 			--14
	if (addfprdy = '1') then state := s15304;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15303; end if;
when s15304 => state := s15305; 	--15
	addfpsclr <= '0';
when s15305 => state := s15306; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15306 => 			--17
	if (addfprdy = '1') then state := s15307;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15306; end if;
when s15307 => state := s15308; 	--18
	addfpsclr <= '0';
when s15308 => state := s15309; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15309 => 			--20
	if (addfprdy = '1') then state := s15310;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15309; end if;
when s15310 => state := s15311; 	--21
	addfpsclr <= '0';
when s15311 => state := s15312; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (751, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15312 => state := s15313; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1440, 12)); -- offset LSB 1392
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s15313 => state := s15314;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1441, 12)); -- offset MSB 1393
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15314 => state := s15315; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15315 => 			--4
	if (fixed2floatrdy = '1') then state := s15316;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15315; end if;
when s15316 => state := s15317; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15317 => 			--6
	if (mulfprdy = '1') then state := s15318;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15317; end if;
when s15318 => state := s15319; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15319 => 			--8
	if (mulfprdy = '1') then state := s15320;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15319; end if;
when s15320 => state := s15321; 	--9
	mulfpsclr <= '0';
when s15321 => state := s15322; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15322 => 			--11
	if (mulfprdy = '1') then state := s15323;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15322; end if;
when s15323 => state := s15324; 	--12
	mulfpsclr <= '0';
when s15324 => state := s15325; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15325 => 			--14
	if (addfprdy = '1') then state := s15326;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15325; end if;
when s15326 => state := s15327; 	--15
	addfpsclr <= '0';
when s15327 => state := s15328; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15328 => 			--17
	if (addfprdy = '1') then state := s15329;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15328; end if;
when s15329 => state := s15330; 	--18
	addfpsclr <= '0';
when s15330 => state := s15331; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15331 => 			--20
	if (addfprdy = '1') then state := s15332;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15331; end if;
when s15332 => state := s15333; 	--21
	addfpsclr <= '0';
when s15333 => state := s15334; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (752, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15334 => state := s15335; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1442, 12)); -- offset LSB 1394
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s15335 => state := s15336;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1443, 12)); -- offset MSB 1395
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15336 => state := s15337; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15337 => 			--4
	if (fixed2floatrdy = '1') then state := s15338;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15337; end if;
when s15338 => state := s15339; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15339 => 			--6
	if (mulfprdy = '1') then state := s15340;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15339; end if;
when s15340 => state := s15341; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15341 => 			--8
	if (mulfprdy = '1') then state := s15342;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15341; end if;
when s15342 => state := s15343; 	--9
	mulfpsclr <= '0';
when s15343 => state := s15344; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15344 => 			--11
	if (mulfprdy = '1') then state := s15345;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15344; end if;
when s15345 => state := s15346; 	--12
	mulfpsclr <= '0';
when s15346 => state := s15347; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15347 => 			--14
	if (addfprdy = '1') then state := s15348;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15347; end if;
when s15348 => state := s15349; 	--15
	addfpsclr <= '0';
when s15349 => state := s15350; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15350 => 			--17
	if (addfprdy = '1') then state := s15351;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15350; end if;
when s15351 => state := s15352; 	--18
	addfpsclr <= '0';
when s15352 => state := s15353; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15353 => 			--20
	if (addfprdy = '1') then state := s15354;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15353; end if;
when s15354 => state := s15355; 	--21
	addfpsclr <= '0';
when s15355 => state := s15356; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (753, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15356 => state := s15357; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1444, 12)); -- offset LSB 1396
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s15357 => state := s15358;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1445, 12)); -- offset MSB 1397
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15358 => state := s15359; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15359 => 			--4
	if (fixed2floatrdy = '1') then state := s15360;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15359; end if;
when s15360 => state := s15361; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15361 => 			--6
	if (mulfprdy = '1') then state := s15362;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15361; end if;
when s15362 => state := s15363; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15363 => 			--8
	if (mulfprdy = '1') then state := s15364;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15363; end if;
when s15364 => state := s15365; 	--9
	mulfpsclr <= '0';
when s15365 => state := s15366; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15366 => 			--11
	if (mulfprdy = '1') then state := s15367;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15366; end if;
when s15367 => state := s15368; 	--12
	mulfpsclr <= '0';
when s15368 => state := s15369; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15369 => 			--14
	if (addfprdy = '1') then state := s15370;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15369; end if;
when s15370 => state := s15371; 	--15
	addfpsclr <= '0';
when s15371 => state := s15372; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15372 => 			--17
	if (addfprdy = '1') then state := s15373;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15372; end if;
when s15373 => state := s15374; 	--18
	addfpsclr <= '0';
when s15374 => state := s15375; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15375 => 			--20
	if (addfprdy = '1') then state := s15376;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15375; end if;
when s15376 => state := s15377; 	--21
	addfpsclr <= '0';
when s15377 => state := s15378; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (754, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15378 => state := s15379; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1446, 12)); -- offset LSB 1398
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s15379 => state := s15380;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1447, 12)); -- offset MSB 1399
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15380 => state := s15381; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15381 => 			--4
	if (fixed2floatrdy = '1') then state := s15382;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15381; end if;
when s15382 => state := s15383; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15383 => 			--6
	if (mulfprdy = '1') then state := s15384;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15383; end if;
when s15384 => state := s15385; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15385 => 			--8
	if (mulfprdy = '1') then state := s15386;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15385; end if;
when s15386 => state := s15387; 	--9
	mulfpsclr <= '0';
when s15387 => state := s15388; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15388 => 			--11
	if (mulfprdy = '1') then state := s15389;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15388; end if;
when s15389 => state := s15390; 	--12
	mulfpsclr <= '0';
when s15390 => state := s15391; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15391 => 			--14
	if (addfprdy = '1') then state := s15392;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15391; end if;
when s15392 => state := s15393; 	--15
	addfpsclr <= '0';
when s15393 => state := s15394; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15394 => 			--17
	if (addfprdy = '1') then state := s15395;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15394; end if;
when s15395 => state := s15396; 	--18
	addfpsclr <= '0';
when s15396 => state := s15397; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15397 => 			--20
	if (addfprdy = '1') then state := s15398;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15397; end if;
when s15398 => state := s15399; 	--21
	addfpsclr <= '0';
when s15399 => state := s15400; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (755, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15400 => state := s15401; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1448, 12)); -- offset LSB 1400
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s15401 => state := s15402;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1449, 12)); -- offset MSB 1401
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15402 => state := s15403; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15403 => 			--4
	if (fixed2floatrdy = '1') then state := s15404;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15403; end if;
when s15404 => state := s15405; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15405 => 			--6
	if (mulfprdy = '1') then state := s15406;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15405; end if;
when s15406 => state := s15407; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15407 => 			--8
	if (mulfprdy = '1') then state := s15408;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15407; end if;
when s15408 => state := s15409; 	--9
	mulfpsclr <= '0';
when s15409 => state := s15410; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15410 => 			--11
	if (mulfprdy = '1') then state := s15411;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15410; end if;
when s15411 => state := s15412; 	--12
	mulfpsclr <= '0';
when s15412 => state := s15413; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15413 => 			--14
	if (addfprdy = '1') then state := s15414;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15413; end if;
when s15414 => state := s15415; 	--15
	addfpsclr <= '0';
when s15415 => state := s15416; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15416 => 			--17
	if (addfprdy = '1') then state := s15417;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15416; end if;
when s15417 => state := s15418; 	--18
	addfpsclr <= '0';
when s15418 => state := s15419; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15419 => 			--20
	if (addfprdy = '1') then state := s15420;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15419; end if;
when s15420 => state := s15421; 	--21
	addfpsclr <= '0';
when s15421 => state := s15422; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (756, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15422 => state := s15423; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1450, 12)); -- offset LSB 1402
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s15423 => state := s15424;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1451, 12)); -- offset MSB 1403
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15424 => state := s15425; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15425 => 			--4
	if (fixed2floatrdy = '1') then state := s15426;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15425; end if;
when s15426 => state := s15427; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15427 => 			--6
	if (mulfprdy = '1') then state := s15428;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15427; end if;
when s15428 => state := s15429; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15429 => 			--8
	if (mulfprdy = '1') then state := s15430;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15429; end if;
when s15430 => state := s15431; 	--9
	mulfpsclr <= '0';
when s15431 => state := s15432; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15432 => 			--11
	if (mulfprdy = '1') then state := s15433;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15432; end if;
when s15433 => state := s15434; 	--12
	mulfpsclr <= '0';
when s15434 => state := s15435; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15435 => 			--14
	if (addfprdy = '1') then state := s15436;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15435; end if;
when s15436 => state := s15437; 	--15
	addfpsclr <= '0';
when s15437 => state := s15438; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15438 => 			--17
	if (addfprdy = '1') then state := s15439;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15438; end if;
when s15439 => state := s15440; 	--18
	addfpsclr <= '0';
when s15440 => state := s15441; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15441 => 			--20
	if (addfprdy = '1') then state := s15442;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15441; end if;
when s15442 => state := s15443; 	--21
	addfpsclr <= '0';
when s15443 => state := s15444; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (757, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15444 => state := s15445; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1452, 12)); -- offset LSB 1404
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s15445 => state := s15446;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1453, 12)); -- offset MSB 1405
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15446 => state := s15447; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15447 => 			--4
	if (fixed2floatrdy = '1') then state := s15448;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15447; end if;
when s15448 => state := s15449; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15449 => 			--6
	if (mulfprdy = '1') then state := s15450;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15449; end if;
when s15450 => state := s15451; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15451 => 			--8
	if (mulfprdy = '1') then state := s15452;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15451; end if;
when s15452 => state := s15453; 	--9
	mulfpsclr <= '0';
when s15453 => state := s15454; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15454 => 			--11
	if (mulfprdy = '1') then state := s15455;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15454; end if;
when s15455 => state := s15456; 	--12
	mulfpsclr <= '0';
when s15456 => state := s15457; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15457 => 			--14
	if (addfprdy = '1') then state := s15458;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15457; end if;
when s15458 => state := s15459; 	--15
	addfpsclr <= '0';
when s15459 => state := s15460; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15460 => 			--17
	if (addfprdy = '1') then state := s15461;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15460; end if;
when s15461 => state := s15462; 	--18
	addfpsclr <= '0';
when s15462 => state := s15463; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15463 => 			--20
	if (addfprdy = '1') then state := s15464;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15463; end if;
when s15464 => state := s15465; 	--21
	addfpsclr <= '0';
when s15465 => state := s15466; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (758, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15466 => state := s15467; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1454, 12)); -- offset LSB 1406
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s15467 => state := s15468;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1455, 12)); -- offset MSB 1407
	addra <= std_logic_vector (to_unsigned (21, 10)); -- OCCrowI 21
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15468 => state := s15469; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15469 => 			--4
	if (fixed2floatrdy = '1') then state := s15470;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15469; end if;
when s15470 => state := s15471; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15471 => 			--6
	if (mulfprdy = '1') then state := s15472;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15471; end if;
when s15472 => state := s15473; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15473 => 			--8
	if (mulfprdy = '1') then state := s15474;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15473; end if;
when s15474 => state := s15475; 	--9
	mulfpsclr <= '0';
when s15475 => state := s15476; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15476 => 			--11
	if (mulfprdy = '1') then state := s15477;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15476; end if;
when s15477 => state := s15478; 	--12
	mulfpsclr <= '0';
when s15478 => state := s15479; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15479 => 			--14
	if (addfprdy = '1') then state := s15480;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15479; end if;
when s15480 => state := s15481; 	--15
	addfpsclr <= '0';
when s15481 => state := s15482; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15482 => 			--17
	if (addfprdy = '1') then state := s15483;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15482; end if;
when s15483 => state := s15484; 	--18
	addfpsclr <= '0';
when s15484 => state := s15485; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15485 => 			--20
	if (addfprdy = '1') then state := s15486;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15485; end if;
when s15486 => state := s15487; 	--21
	addfpsclr <= '0';
when s15487 => state := s15488; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (759, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15488 => state := s15489; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1456, 12)); -- offset LSB 1408
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s15489 => state := s15490;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1457, 12)); -- offset MSB 1409
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15490 => state := s15491; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15491 => 			--4
	if (fixed2floatrdy = '1') then state := s15492;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15491; end if;
when s15492 => state := s15493; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15493 => 			--6
	if (mulfprdy = '1') then state := s15494;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15493; end if;
when s15494 => state := s15495; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15495 => 			--8
	if (mulfprdy = '1') then state := s15496;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15495; end if;
when s15496 => state := s15497; 	--9
	mulfpsclr <= '0';
when s15497 => state := s15498; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15498 => 			--11
	if (mulfprdy = '1') then state := s15499;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15498; end if;
when s15499 => state := s15500; 	--12
	mulfpsclr <= '0';
when s15500 => state := s15501; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15501 => 			--14
	if (addfprdy = '1') then state := s15502;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15501; end if;
when s15502 => state := s15503; 	--15
	addfpsclr <= '0';
when s15503 => state := s15504; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15504 => 			--17
	if (addfprdy = '1') then state := s15505;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15504; end if;
when s15505 => state := s15506; 	--18
	addfpsclr <= '0';
when s15506 => state := s15507; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15507 => 			--20
	if (addfprdy = '1') then state := s15508;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15507; end if;
when s15508 => state := s15509; 	--21
	addfpsclr <= '0';
when s15509 => state := s15510; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (760, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15510 => state := s15511; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1458, 12)); -- offset LSB 1410
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s15511 => state := s15512;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1459, 12)); -- offset MSB 1411
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15512 => state := s15513; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15513 => 			--4
	if (fixed2floatrdy = '1') then state := s15514;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15513; end if;
when s15514 => state := s15515; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15515 => 			--6
	if (mulfprdy = '1') then state := s15516;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15515; end if;
when s15516 => state := s15517; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15517 => 			--8
	if (mulfprdy = '1') then state := s15518;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15517; end if;
when s15518 => state := s15519; 	--9
	mulfpsclr <= '0';
when s15519 => state := s15520; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15520 => 			--11
	if (mulfprdy = '1') then state := s15521;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15520; end if;
when s15521 => state := s15522; 	--12
	mulfpsclr <= '0';
when s15522 => state := s15523; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15523 => 			--14
	if (addfprdy = '1') then state := s15524;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15523; end if;
when s15524 => state := s15525; 	--15
	addfpsclr <= '0';
when s15525 => state := s15526; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15526 => 			--17
	if (addfprdy = '1') then state := s15527;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15526; end if;
when s15527 => state := s15528; 	--18
	addfpsclr <= '0';
when s15528 => state := s15529; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15529 => 			--20
	if (addfprdy = '1') then state := s15530;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15529; end if;
when s15530 => state := s15531; 	--21
	addfpsclr <= '0';
when s15531 => state := s15532; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (761, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15532 => state := s15533; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1460, 12)); -- offset LSB 1412
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s15533 => state := s15534;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1461, 12)); -- offset MSB 1413
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15534 => state := s15535; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15535 => 			--4
	if (fixed2floatrdy = '1') then state := s15536;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15535; end if;
when s15536 => state := s15537; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15537 => 			--6
	if (mulfprdy = '1') then state := s15538;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15537; end if;
when s15538 => state := s15539; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15539 => 			--8
	if (mulfprdy = '1') then state := s15540;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15539; end if;
when s15540 => state := s15541; 	--9
	mulfpsclr <= '0';
when s15541 => state := s15542; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15542 => 			--11
	if (mulfprdy = '1') then state := s15543;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15542; end if;
when s15543 => state := s15544; 	--12
	mulfpsclr <= '0';
when s15544 => state := s15545; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15545 => 			--14
	if (addfprdy = '1') then state := s15546;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15545; end if;
when s15546 => state := s15547; 	--15
	addfpsclr <= '0';
when s15547 => state := s15548; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15548 => 			--17
	if (addfprdy = '1') then state := s15549;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15548; end if;
when s15549 => state := s15550; 	--18
	addfpsclr <= '0';
when s15550 => state := s15551; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15551 => 			--20
	if (addfprdy = '1') then state := s15552;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15551; end if;
when s15552 => state := s15553; 	--21
	addfpsclr <= '0';
when s15553 => state := s15554; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (762, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15554 => state := s15555; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1462, 12)); -- offset LSB 1414
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s15555 => state := s15556;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1463, 12)); -- offset MSB 1415
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15556 => state := s15557; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15557 => 			--4
	if (fixed2floatrdy = '1') then state := s15558;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15557; end if;
when s15558 => state := s15559; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15559 => 			--6
	if (mulfprdy = '1') then state := s15560;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15559; end if;
when s15560 => state := s15561; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15561 => 			--8
	if (mulfprdy = '1') then state := s15562;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15561; end if;
when s15562 => state := s15563; 	--9
	mulfpsclr <= '0';
when s15563 => state := s15564; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15564 => 			--11
	if (mulfprdy = '1') then state := s15565;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15564; end if;
when s15565 => state := s15566; 	--12
	mulfpsclr <= '0';
when s15566 => state := s15567; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15567 => 			--14
	if (addfprdy = '1') then state := s15568;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15567; end if;
when s15568 => state := s15569; 	--15
	addfpsclr <= '0';
when s15569 => state := s15570; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15570 => 			--17
	if (addfprdy = '1') then state := s15571;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15570; end if;
when s15571 => state := s15572; 	--18
	addfpsclr <= '0';
when s15572 => state := s15573; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15573 => 			--20
	if (addfprdy = '1') then state := s15574;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15573; end if;
when s15574 => state := s15575; 	--21
	addfpsclr <= '0';
when s15575 => state := s15576; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (763, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15576 => state := s15577; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1464, 12)); -- offset LSB 1416
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s15577 => state := s15578;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1465, 12)); -- offset MSB 1417
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15578 => state := s15579; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15579 => 			--4
	if (fixed2floatrdy = '1') then state := s15580;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15579; end if;
when s15580 => state := s15581; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15581 => 			--6
	if (mulfprdy = '1') then state := s15582;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15581; end if;
when s15582 => state := s15583; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15583 => 			--8
	if (mulfprdy = '1') then state := s15584;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15583; end if;
when s15584 => state := s15585; 	--9
	mulfpsclr <= '0';
when s15585 => state := s15586; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15586 => 			--11
	if (mulfprdy = '1') then state := s15587;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15586; end if;
when s15587 => state := s15588; 	--12
	mulfpsclr <= '0';
when s15588 => state := s15589; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15589 => 			--14
	if (addfprdy = '1') then state := s15590;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15589; end if;
when s15590 => state := s15591; 	--15
	addfpsclr <= '0';
when s15591 => state := s15592; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15592 => 			--17
	if (addfprdy = '1') then state := s15593;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15592; end if;
when s15593 => state := s15594; 	--18
	addfpsclr <= '0';
when s15594 => state := s15595; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15595 => 			--20
	if (addfprdy = '1') then state := s15596;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15595; end if;
when s15596 => state := s15597; 	--21
	addfpsclr <= '0';
when s15597 => state := s15598; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (764, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15598 => state := s15599; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1466, 12)); -- offset LSB 1418
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s15599 => state := s15600;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1467, 12)); -- offset MSB 1419
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15600 => state := s15601; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15601 => 			--4
	if (fixed2floatrdy = '1') then state := s15602;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15601; end if;
when s15602 => state := s15603; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15603 => 			--6
	if (mulfprdy = '1') then state := s15604;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15603; end if;
when s15604 => state := s15605; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15605 => 			--8
	if (mulfprdy = '1') then state := s15606;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15605; end if;
when s15606 => state := s15607; 	--9
	mulfpsclr <= '0';
when s15607 => state := s15608; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15608 => 			--11
	if (mulfprdy = '1') then state := s15609;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15608; end if;
when s15609 => state := s15610; 	--12
	mulfpsclr <= '0';
when s15610 => state := s15611; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15611 => 			--14
	if (addfprdy = '1') then state := s15612;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15611; end if;
when s15612 => state := s15613; 	--15
	addfpsclr <= '0';
when s15613 => state := s15614; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15614 => 			--17
	if (addfprdy = '1') then state := s15615;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15614; end if;
when s15615 => state := s15616; 	--18
	addfpsclr <= '0';
when s15616 => state := s15617; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15617 => 			--20
	if (addfprdy = '1') then state := s15618;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15617; end if;
when s15618 => state := s15619; 	--21
	addfpsclr <= '0';
when s15619 => state := s15620; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (765, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15620 => state := s15621; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1468, 12)); -- offset LSB 1420
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s15621 => state := s15622;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1469, 12)); -- offset MSB 1421
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15622 => state := s15623; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15623 => 			--4
	if (fixed2floatrdy = '1') then state := s15624;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15623; end if;
when s15624 => state := s15625; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15625 => 			--6
	if (mulfprdy = '1') then state := s15626;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15625; end if;
when s15626 => state := s15627; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15627 => 			--8
	if (mulfprdy = '1') then state := s15628;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15627; end if;
when s15628 => state := s15629; 	--9
	mulfpsclr <= '0';
when s15629 => state := s15630; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15630 => 			--11
	if (mulfprdy = '1') then state := s15631;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15630; end if;
when s15631 => state := s15632; 	--12
	mulfpsclr <= '0';
when s15632 => state := s15633; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15633 => 			--14
	if (addfprdy = '1') then state := s15634;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15633; end if;
when s15634 => state := s15635; 	--15
	addfpsclr <= '0';
when s15635 => state := s15636; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15636 => 			--17
	if (addfprdy = '1') then state := s15637;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15636; end if;
when s15637 => state := s15638; 	--18
	addfpsclr <= '0';
when s15638 => state := s15639; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15639 => 			--20
	if (addfprdy = '1') then state := s15640;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15639; end if;
when s15640 => state := s15641; 	--21
	addfpsclr <= '0';
when s15641 => state := s15642; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (766, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15642 => state := s15643; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1470, 12)); -- offset LSB 1422
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s15643 => state := s15644;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1471, 12)); -- offset MSB 1423
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15644 => state := s15645; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15645 => 			--4
	if (fixed2floatrdy = '1') then state := s15646;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15645; end if;
when s15646 => state := s15647; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15647 => 			--6
	if (mulfprdy = '1') then state := s15648;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15647; end if;
when s15648 => state := s15649; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15649 => 			--8
	if (mulfprdy = '1') then state := s15650;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15649; end if;
when s15650 => state := s15651; 	--9
	mulfpsclr <= '0';
when s15651 => state := s15652; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15652 => 			--11
	if (mulfprdy = '1') then state := s15653;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15652; end if;
when s15653 => state := s15654; 	--12
	mulfpsclr <= '0';
when s15654 => state := s15655; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15655 => 			--14
	if (addfprdy = '1') then state := s15656;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15655; end if;
when s15656 => state := s15657; 	--15
	addfpsclr <= '0';
when s15657 => state := s15658; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15658 => 			--17
	if (addfprdy = '1') then state := s15659;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15658; end if;
when s15659 => state := s15660; 	--18
	addfpsclr <= '0';
when s15660 => state := s15661; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15661 => 			--20
	if (addfprdy = '1') then state := s15662;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15661; end if;
when s15662 => state := s15663; 	--21
	addfpsclr <= '0';
when s15663 => state := s15664; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (767, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15664 => state := s15665; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1472, 12)); -- offset LSB 1424
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s15665 => state := s15666;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1473, 12)); -- offset MSB 1425
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15666 => state := s15667; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15667 => 			--4
	if (fixed2floatrdy = '1') then state := s15668;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15667; end if;
when s15668 => state := s15669; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15669 => 			--6
	if (mulfprdy = '1') then state := s15670;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15669; end if;
when s15670 => state := s15671; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15671 => 			--8
	if (mulfprdy = '1') then state := s15672;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15671; end if;
when s15672 => state := s15673; 	--9
	mulfpsclr <= '0';
when s15673 => state := s15674; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15674 => 			--11
	if (mulfprdy = '1') then state := s15675;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15674; end if;
when s15675 => state := s15676; 	--12
	mulfpsclr <= '0';
when s15676 => state := s15677; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15677 => 			--14
	if (addfprdy = '1') then state := s15678;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15677; end if;
when s15678 => state := s15679; 	--15
	addfpsclr <= '0';
when s15679 => state := s15680; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15680 => 			--17
	if (addfprdy = '1') then state := s15681;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15680; end if;
when s15681 => state := s15682; 	--18
	addfpsclr <= '0';
when s15682 => state := s15683; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15683 => 			--20
	if (addfprdy = '1') then state := s15684;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15683; end if;
when s15684 => state := s15685; 	--21
	addfpsclr <= '0';
when s15685 => state := s15686; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (768, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15686 => state := s15687; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1474, 12)); -- offset LSB 1426
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s15687 => state := s15688;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1475, 12)); -- offset MSB 1427
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15688 => state := s15689; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15689 => 			--4
	if (fixed2floatrdy = '1') then state := s15690;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15689; end if;
when s15690 => state := s15691; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15691 => 			--6
	if (mulfprdy = '1') then state := s15692;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15691; end if;
when s15692 => state := s15693; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15693 => 			--8
	if (mulfprdy = '1') then state := s15694;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15693; end if;
when s15694 => state := s15695; 	--9
	mulfpsclr <= '0';
when s15695 => state := s15696; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15696 => 			--11
	if (mulfprdy = '1') then state := s15697;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15696; end if;
when s15697 => state := s15698; 	--12
	mulfpsclr <= '0';
when s15698 => state := s15699; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15699 => 			--14
	if (addfprdy = '1') then state := s15700;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15699; end if;
when s15700 => state := s15701; 	--15
	addfpsclr <= '0';
when s15701 => state := s15702; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15702 => 			--17
	if (addfprdy = '1') then state := s15703;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15702; end if;
when s15703 => state := s15704; 	--18
	addfpsclr <= '0';
when s15704 => state := s15705; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15705 => 			--20
	if (addfprdy = '1') then state := s15706;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15705; end if;
when s15706 => state := s15707; 	--21
	addfpsclr <= '0';
when s15707 => state := s15708; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (769, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15708 => state := s15709; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1476, 12)); -- offset LSB 1428
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s15709 => state := s15710;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1477, 12)); -- offset MSB 1429
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15710 => state := s15711; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15711 => 			--4
	if (fixed2floatrdy = '1') then state := s15712;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15711; end if;
when s15712 => state := s15713; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15713 => 			--6
	if (mulfprdy = '1') then state := s15714;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15713; end if;
when s15714 => state := s15715; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15715 => 			--8
	if (mulfprdy = '1') then state := s15716;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15715; end if;
when s15716 => state := s15717; 	--9
	mulfpsclr <= '0';
when s15717 => state := s15718; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15718 => 			--11
	if (mulfprdy = '1') then state := s15719;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15718; end if;
when s15719 => state := s15720; 	--12
	mulfpsclr <= '0';
when s15720 => state := s15721; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15721 => 			--14
	if (addfprdy = '1') then state := s15722;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15721; end if;
when s15722 => state := s15723; 	--15
	addfpsclr <= '0';
when s15723 => state := s15724; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15724 => 			--17
	if (addfprdy = '1') then state := s15725;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15724; end if;
when s15725 => state := s15726; 	--18
	addfpsclr <= '0';
when s15726 => state := s15727; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15727 => 			--20
	if (addfprdy = '1') then state := s15728;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15727; end if;
when s15728 => state := s15729; 	--21
	addfpsclr <= '0';
when s15729 => state := s15730; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (770, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15730 => state := s15731; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1478, 12)); -- offset LSB 1430
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s15731 => state := s15732;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1479, 12)); -- offset MSB 1431
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15732 => state := s15733; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15733 => 			--4
	if (fixed2floatrdy = '1') then state := s15734;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15733; end if;
when s15734 => state := s15735; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15735 => 			--6
	if (mulfprdy = '1') then state := s15736;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15735; end if;
when s15736 => state := s15737; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15737 => 			--8
	if (mulfprdy = '1') then state := s15738;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15737; end if;
when s15738 => state := s15739; 	--9
	mulfpsclr <= '0';
when s15739 => state := s15740; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15740 => 			--11
	if (mulfprdy = '1') then state := s15741;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15740; end if;
when s15741 => state := s15742; 	--12
	mulfpsclr <= '0';
when s15742 => state := s15743; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15743 => 			--14
	if (addfprdy = '1') then state := s15744;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15743; end if;
when s15744 => state := s15745; 	--15
	addfpsclr <= '0';
when s15745 => state := s15746; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15746 => 			--17
	if (addfprdy = '1') then state := s15747;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15746; end if;
when s15747 => state := s15748; 	--18
	addfpsclr <= '0';
when s15748 => state := s15749; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15749 => 			--20
	if (addfprdy = '1') then state := s15750;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15749; end if;
when s15750 => state := s15751; 	--21
	addfpsclr <= '0';
when s15751 => state := s15752; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (771, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15752 => state := s15753; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1480, 12)); -- offset LSB 1432
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s15753 => state := s15754;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1481, 12)); -- offset MSB 1433
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15754 => state := s15755; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15755 => 			--4
	if (fixed2floatrdy = '1') then state := s15756;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15755; end if;
when s15756 => state := s15757; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15757 => 			--6
	if (mulfprdy = '1') then state := s15758;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15757; end if;
when s15758 => state := s15759; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15759 => 			--8
	if (mulfprdy = '1') then state := s15760;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15759; end if;
when s15760 => state := s15761; 	--9
	mulfpsclr <= '0';
when s15761 => state := s15762; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15762 => 			--11
	if (mulfprdy = '1') then state := s15763;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15762; end if;
when s15763 => state := s15764; 	--12
	mulfpsclr <= '0';
when s15764 => state := s15765; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15765 => 			--14
	if (addfprdy = '1') then state := s15766;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15765; end if;
when s15766 => state := s15767; 	--15
	addfpsclr <= '0';
when s15767 => state := s15768; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15768 => 			--17
	if (addfprdy = '1') then state := s15769;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15768; end if;
when s15769 => state := s15770; 	--18
	addfpsclr <= '0';
when s15770 => state := s15771; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15771 => 			--20
	if (addfprdy = '1') then state := s15772;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15771; end if;
when s15772 => state := s15773; 	--21
	addfpsclr <= '0';
when s15773 => state := s15774; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (772, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15774 => state := s15775; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1482, 12)); -- offset LSB 1434
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s15775 => state := s15776;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1483, 12)); -- offset MSB 1435
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15776 => state := s15777; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15777 => 			--4
	if (fixed2floatrdy = '1') then state := s15778;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15777; end if;
when s15778 => state := s15779; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15779 => 			--6
	if (mulfprdy = '1') then state := s15780;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15779; end if;
when s15780 => state := s15781; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15781 => 			--8
	if (mulfprdy = '1') then state := s15782;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15781; end if;
when s15782 => state := s15783; 	--9
	mulfpsclr <= '0';
when s15783 => state := s15784; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15784 => 			--11
	if (mulfprdy = '1') then state := s15785;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15784; end if;
when s15785 => state := s15786; 	--12
	mulfpsclr <= '0';
when s15786 => state := s15787; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15787 => 			--14
	if (addfprdy = '1') then state := s15788;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15787; end if;
when s15788 => state := s15789; 	--15
	addfpsclr <= '0';
when s15789 => state := s15790; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15790 => 			--17
	if (addfprdy = '1') then state := s15791;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15790; end if;
when s15791 => state := s15792; 	--18
	addfpsclr <= '0';
when s15792 => state := s15793; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15793 => 			--20
	if (addfprdy = '1') then state := s15794;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15793; end if;
when s15794 => state := s15795; 	--21
	addfpsclr <= '0';
when s15795 => state := s15796; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (773, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15796 => state := s15797; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1484, 12)); -- offset LSB 1436
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s15797 => state := s15798;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1485, 12)); -- offset MSB 1437
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15798 => state := s15799; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15799 => 			--4
	if (fixed2floatrdy = '1') then state := s15800;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15799; end if;
when s15800 => state := s15801; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15801 => 			--6
	if (mulfprdy = '1') then state := s15802;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15801; end if;
when s15802 => state := s15803; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15803 => 			--8
	if (mulfprdy = '1') then state := s15804;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15803; end if;
when s15804 => state := s15805; 	--9
	mulfpsclr <= '0';
when s15805 => state := s15806; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15806 => 			--11
	if (mulfprdy = '1') then state := s15807;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15806; end if;
when s15807 => state := s15808; 	--12
	mulfpsclr <= '0';
when s15808 => state := s15809; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15809 => 			--14
	if (addfprdy = '1') then state := s15810;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15809; end if;
when s15810 => state := s15811; 	--15
	addfpsclr <= '0';
when s15811 => state := s15812; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15812 => 			--17
	if (addfprdy = '1') then state := s15813;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15812; end if;
when s15813 => state := s15814; 	--18
	addfpsclr <= '0';
when s15814 => state := s15815; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15815 => 			--20
	if (addfprdy = '1') then state := s15816;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15815; end if;
when s15816 => state := s15817; 	--21
	addfpsclr <= '0';
when s15817 => state := s15818; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (774, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15818 => state := s15819; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1486, 12)); -- offset LSB 1438
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s15819 => state := s15820;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1487, 12)); -- offset MSB 1439
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15820 => state := s15821; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15821 => 			--4
	if (fixed2floatrdy = '1') then state := s15822;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15821; end if;
when s15822 => state := s15823; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15823 => 			--6
	if (mulfprdy = '1') then state := s15824;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15823; end if;
when s15824 => state := s15825; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15825 => 			--8
	if (mulfprdy = '1') then state := s15826;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15825; end if;
when s15826 => state := s15827; 	--9
	mulfpsclr <= '0';
when s15827 => state := s15828; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15828 => 			--11
	if (mulfprdy = '1') then state := s15829;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15828; end if;
when s15829 => state := s15830; 	--12
	mulfpsclr <= '0';
when s15830 => state := s15831; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15831 => 			--14
	if (addfprdy = '1') then state := s15832;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15831; end if;
when s15832 => state := s15833; 	--15
	addfpsclr <= '0';
when s15833 => state := s15834; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15834 => 			--17
	if (addfprdy = '1') then state := s15835;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15834; end if;
when s15835 => state := s15836; 	--18
	addfpsclr <= '0';
when s15836 => state := s15837; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15837 => 			--20
	if (addfprdy = '1') then state := s15838;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15837; end if;
when s15838 => state := s15839; 	--21
	addfpsclr <= '0';
when s15839 => state := s15840; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (775, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15840 => state := s15841; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1488, 12)); -- offset LSB 1440
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s15841 => state := s15842;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1489, 12)); -- offset MSB 1441
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15842 => state := s15843; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15843 => 			--4
	if (fixed2floatrdy = '1') then state := s15844;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15843; end if;
when s15844 => state := s15845; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15845 => 			--6
	if (mulfprdy = '1') then state := s15846;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15845; end if;
when s15846 => state := s15847; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15847 => 			--8
	if (mulfprdy = '1') then state := s15848;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15847; end if;
when s15848 => state := s15849; 	--9
	mulfpsclr <= '0';
when s15849 => state := s15850; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15850 => 			--11
	if (mulfprdy = '1') then state := s15851;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15850; end if;
when s15851 => state := s15852; 	--12
	mulfpsclr <= '0';
when s15852 => state := s15853; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15853 => 			--14
	if (addfprdy = '1') then state := s15854;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15853; end if;
when s15854 => state := s15855; 	--15
	addfpsclr <= '0';
when s15855 => state := s15856; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15856 => 			--17
	if (addfprdy = '1') then state := s15857;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15856; end if;
when s15857 => state := s15858; 	--18
	addfpsclr <= '0';
when s15858 => state := s15859; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15859 => 			--20
	if (addfprdy = '1') then state := s15860;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15859; end if;
when s15860 => state := s15861; 	--21
	addfpsclr <= '0';
when s15861 => state := s15862; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (776, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15862 => state := s15863; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1490, 12)); -- offset LSB 1442
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s15863 => state := s15864;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1491, 12)); -- offset MSB 1443
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15864 => state := s15865; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15865 => 			--4
	if (fixed2floatrdy = '1') then state := s15866;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15865; end if;
when s15866 => state := s15867; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15867 => 			--6
	if (mulfprdy = '1') then state := s15868;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15867; end if;
when s15868 => state := s15869; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15869 => 			--8
	if (mulfprdy = '1') then state := s15870;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15869; end if;
when s15870 => state := s15871; 	--9
	mulfpsclr <= '0';
when s15871 => state := s15872; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15872 => 			--11
	if (mulfprdy = '1') then state := s15873;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15872; end if;
when s15873 => state := s15874; 	--12
	mulfpsclr <= '0';
when s15874 => state := s15875; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15875 => 			--14
	if (addfprdy = '1') then state := s15876;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15875; end if;
when s15876 => state := s15877; 	--15
	addfpsclr <= '0';
when s15877 => state := s15878; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15878 => 			--17
	if (addfprdy = '1') then state := s15879;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15878; end if;
when s15879 => state := s15880; 	--18
	addfpsclr <= '0';
when s15880 => state := s15881; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15881 => 			--20
	if (addfprdy = '1') then state := s15882;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15881; end if;
when s15882 => state := s15883; 	--21
	addfpsclr <= '0';
when s15883 => state := s15884; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (777, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15884 => state := s15885; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1492, 12)); -- offset LSB 1444
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s15885 => state := s15886;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1493, 12)); -- offset MSB 1445
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15886 => state := s15887; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15887 => 			--4
	if (fixed2floatrdy = '1') then state := s15888;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15887; end if;
when s15888 => state := s15889; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15889 => 			--6
	if (mulfprdy = '1') then state := s15890;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15889; end if;
when s15890 => state := s15891; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15891 => 			--8
	if (mulfprdy = '1') then state := s15892;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15891; end if;
when s15892 => state := s15893; 	--9
	mulfpsclr <= '0';
when s15893 => state := s15894; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15894 => 			--11
	if (mulfprdy = '1') then state := s15895;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15894; end if;
when s15895 => state := s15896; 	--12
	mulfpsclr <= '0';
when s15896 => state := s15897; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15897 => 			--14
	if (addfprdy = '1') then state := s15898;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15897; end if;
when s15898 => state := s15899; 	--15
	addfpsclr <= '0';
when s15899 => state := s15900; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15900 => 			--17
	if (addfprdy = '1') then state := s15901;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15900; end if;
when s15901 => state := s15902; 	--18
	addfpsclr <= '0';
when s15902 => state := s15903; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15903 => 			--20
	if (addfprdy = '1') then state := s15904;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15903; end if;
when s15904 => state := s15905; 	--21
	addfpsclr <= '0';
when s15905 => state := s15906; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (778, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15906 => state := s15907; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1494, 12)); -- offset LSB 1446
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s15907 => state := s15908;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1495, 12)); -- offset MSB 1447
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15908 => state := s15909; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15909 => 			--4
	if (fixed2floatrdy = '1') then state := s15910;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15909; end if;
when s15910 => state := s15911; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15911 => 			--6
	if (mulfprdy = '1') then state := s15912;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15911; end if;
when s15912 => state := s15913; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15913 => 			--8
	if (mulfprdy = '1') then state := s15914;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15913; end if;
when s15914 => state := s15915; 	--9
	mulfpsclr <= '0';
when s15915 => state := s15916; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15916 => 			--11
	if (mulfprdy = '1') then state := s15917;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15916; end if;
when s15917 => state := s15918; 	--12
	mulfpsclr <= '0';
when s15918 => state := s15919; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15919 => 			--14
	if (addfprdy = '1') then state := s15920;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15919; end if;
when s15920 => state := s15921; 	--15
	addfpsclr <= '0';
when s15921 => state := s15922; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15922 => 			--17
	if (addfprdy = '1') then state := s15923;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15922; end if;
when s15923 => state := s15924; 	--18
	addfpsclr <= '0';
when s15924 => state := s15925; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15925 => 			--20
	if (addfprdy = '1') then state := s15926;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15925; end if;
when s15926 => state := s15927; 	--21
	addfpsclr <= '0';
when s15927 => state := s15928; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (779, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15928 => state := s15929; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1496, 12)); -- offset LSB 1448
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s15929 => state := s15930;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1497, 12)); -- offset MSB 1449
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15930 => state := s15931; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15931 => 			--4
	if (fixed2floatrdy = '1') then state := s15932;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15931; end if;
when s15932 => state := s15933; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15933 => 			--6
	if (mulfprdy = '1') then state := s15934;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15933; end if;
when s15934 => state := s15935; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15935 => 			--8
	if (mulfprdy = '1') then state := s15936;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15935; end if;
when s15936 => state := s15937; 	--9
	mulfpsclr <= '0';
when s15937 => state := s15938; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15938 => 			--11
	if (mulfprdy = '1') then state := s15939;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15938; end if;
when s15939 => state := s15940; 	--12
	mulfpsclr <= '0';
when s15940 => state := s15941; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15941 => 			--14
	if (addfprdy = '1') then state := s15942;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15941; end if;
when s15942 => state := s15943; 	--15
	addfpsclr <= '0';
when s15943 => state := s15944; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15944 => 			--17
	if (addfprdy = '1') then state := s15945;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15944; end if;
when s15945 => state := s15946; 	--18
	addfpsclr <= '0';
when s15946 => state := s15947; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15947 => 			--20
	if (addfprdy = '1') then state := s15948;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15947; end if;
when s15948 => state := s15949; 	--21
	addfpsclr <= '0';
when s15949 => state := s15950; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (780, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15950 => state := s15951; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1498, 12)); -- offset LSB 1450
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s15951 => state := s15952;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1499, 12)); -- offset MSB 1451
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15952 => state := s15953; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15953 => 			--4
	if (fixed2floatrdy = '1') then state := s15954;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15953; end if;
when s15954 => state := s15955; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15955 => 			--6
	if (mulfprdy = '1') then state := s15956;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15955; end if;
when s15956 => state := s15957; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15957 => 			--8
	if (mulfprdy = '1') then state := s15958;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15957; end if;
when s15958 => state := s15959; 	--9
	mulfpsclr <= '0';
when s15959 => state := s15960; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15960 => 			--11
	if (mulfprdy = '1') then state := s15961;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15960; end if;
when s15961 => state := s15962; 	--12
	mulfpsclr <= '0';
when s15962 => state := s15963; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15963 => 			--14
	if (addfprdy = '1') then state := s15964;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15963; end if;
when s15964 => state := s15965; 	--15
	addfpsclr <= '0';
when s15965 => state := s15966; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15966 => 			--17
	if (addfprdy = '1') then state := s15967;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15966; end if;
when s15967 => state := s15968; 	--18
	addfpsclr <= '0';
when s15968 => state := s15969; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15969 => 			--20
	if (addfprdy = '1') then state := s15970;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15969; end if;
when s15970 => state := s15971; 	--21
	addfpsclr <= '0';
when s15971 => state := s15972; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (781, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15972 => state := s15973; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1500, 12)); -- offset LSB 1452
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s15973 => state := s15974;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1501, 12)); -- offset MSB 1453
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15974 => state := s15975; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15975 => 			--4
	if (fixed2floatrdy = '1') then state := s15976;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15975; end if;
when s15976 => state := s15977; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15977 => 			--6
	if (mulfprdy = '1') then state := s15978;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15977; end if;
when s15978 => state := s15979; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s15979 => 			--8
	if (mulfprdy = '1') then state := s15980;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15979; end if;
when s15980 => state := s15981; 	--9
	mulfpsclr <= '0';
when s15981 => state := s15982; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s15982 => 			--11
	if (mulfprdy = '1') then state := s15983;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15982; end if;
when s15983 => state := s15984; 	--12
	mulfpsclr <= '0';
when s15984 => state := s15985; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s15985 => 			--14
	if (addfprdy = '1') then state := s15986;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15985; end if;
when s15986 => state := s15987; 	--15
	addfpsclr <= '0';
when s15987 => state := s15988; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s15988 => 			--17
	if (addfprdy = '1') then state := s15989;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15988; end if;
when s15989 => state := s15990; 	--18
	addfpsclr <= '0';
when s15990 => state := s15991; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s15991 => 			--20
	if (addfprdy = '1') then state := s15992;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s15991; end if;
when s15992 => state := s15993; 	--21
	addfpsclr <= '0';
when s15993 => state := s15994; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (782, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s15994 => state := s15995; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1502, 12)); -- offset LSB 1454
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s15995 => state := s15996;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1503, 12)); -- offset MSB 1455
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s15996 => state := s15997; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s15997 => 			--4
	if (fixed2floatrdy = '1') then state := s15998;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s15997; end if;
when s15998 => state := s15999; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s15999 => 			--6
	if (mulfprdy = '1') then state := s16000;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s15999; end if;
when s16000 => state := s16001; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16001 => 			--8
	if (mulfprdy = '1') then state := s16002;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16001; end if;
when s16002 => state := s16003; 	--9
	mulfpsclr <= '0';
when s16003 => state := s16004; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16004 => 			--11
	if (mulfprdy = '1') then state := s16005;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16004; end if;
when s16005 => state := s16006; 	--12
	mulfpsclr <= '0';
when s16006 => state := s16007; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16007 => 			--14
	if (addfprdy = '1') then state := s16008;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16007; end if;
when s16008 => state := s16009; 	--15
	addfpsclr <= '0';
when s16009 => state := s16010; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16010 => 			--17
	if (addfprdy = '1') then state := s16011;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16010; end if;
when s16011 => state := s16012; 	--18
	addfpsclr <= '0';
when s16012 => state := s16013; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16013 => 			--20
	if (addfprdy = '1') then state := s16014;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16013; end if;
when s16014 => state := s16015; 	--21
	addfpsclr <= '0';
when s16015 => state := s16016; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (783, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16016 => state := s16017; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1504, 12)); -- offset LSB 1456
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s16017 => state := s16018;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1505, 12)); -- offset MSB 1457
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16018 => state := s16019; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16019 => 			--4
	if (fixed2floatrdy = '1') then state := s16020;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16019; end if;
when s16020 => state := s16021; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16021 => 			--6
	if (mulfprdy = '1') then state := s16022;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16021; end if;
when s16022 => state := s16023; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16023 => 			--8
	if (mulfprdy = '1') then state := s16024;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16023; end if;
when s16024 => state := s16025; 	--9
	mulfpsclr <= '0';
when s16025 => state := s16026; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16026 => 			--11
	if (mulfprdy = '1') then state := s16027;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16026; end if;
when s16027 => state := s16028; 	--12
	mulfpsclr <= '0';
when s16028 => state := s16029; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16029 => 			--14
	if (addfprdy = '1') then state := s16030;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16029; end if;
when s16030 => state := s16031; 	--15
	addfpsclr <= '0';
when s16031 => state := s16032; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16032 => 			--17
	if (addfprdy = '1') then state := s16033;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16032; end if;
when s16033 => state := s16034; 	--18
	addfpsclr <= '0';
when s16034 => state := s16035; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16035 => 			--20
	if (addfprdy = '1') then state := s16036;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16035; end if;
when s16036 => state := s16037; 	--21
	addfpsclr <= '0';
when s16037 => state := s16038; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (784, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16038 => state := s16039; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1506, 12)); -- offset LSB 1458
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s16039 => state := s16040;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1507, 12)); -- offset MSB 1459
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16040 => state := s16041; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16041 => 			--4
	if (fixed2floatrdy = '1') then state := s16042;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16041; end if;
when s16042 => state := s16043; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16043 => 			--6
	if (mulfprdy = '1') then state := s16044;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16043; end if;
when s16044 => state := s16045; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16045 => 			--8
	if (mulfprdy = '1') then state := s16046;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16045; end if;
when s16046 => state := s16047; 	--9
	mulfpsclr <= '0';
when s16047 => state := s16048; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16048 => 			--11
	if (mulfprdy = '1') then state := s16049;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16048; end if;
when s16049 => state := s16050; 	--12
	mulfpsclr <= '0';
when s16050 => state := s16051; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16051 => 			--14
	if (addfprdy = '1') then state := s16052;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16051; end if;
when s16052 => state := s16053; 	--15
	addfpsclr <= '0';
when s16053 => state := s16054; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16054 => 			--17
	if (addfprdy = '1') then state := s16055;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16054; end if;
when s16055 => state := s16056; 	--18
	addfpsclr <= '0';
when s16056 => state := s16057; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16057 => 			--20
	if (addfprdy = '1') then state := s16058;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16057; end if;
when s16058 => state := s16059; 	--21
	addfpsclr <= '0';
when s16059 => state := s16060; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (785, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16060 => state := s16061; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1508, 12)); -- offset LSB 1460
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s16061 => state := s16062;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1509, 12)); -- offset MSB 1461
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16062 => state := s16063; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16063 => 			--4
	if (fixed2floatrdy = '1') then state := s16064;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16063; end if;
when s16064 => state := s16065; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16065 => 			--6
	if (mulfprdy = '1') then state := s16066;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16065; end if;
when s16066 => state := s16067; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16067 => 			--8
	if (mulfprdy = '1') then state := s16068;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16067; end if;
when s16068 => state := s16069; 	--9
	mulfpsclr <= '0';
when s16069 => state := s16070; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16070 => 			--11
	if (mulfprdy = '1') then state := s16071;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16070; end if;
when s16071 => state := s16072; 	--12
	mulfpsclr <= '0';
when s16072 => state := s16073; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16073 => 			--14
	if (addfprdy = '1') then state := s16074;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16073; end if;
when s16074 => state := s16075; 	--15
	addfpsclr <= '0';
when s16075 => state := s16076; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16076 => 			--17
	if (addfprdy = '1') then state := s16077;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16076; end if;
when s16077 => state := s16078; 	--18
	addfpsclr <= '0';
when s16078 => state := s16079; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16079 => 			--20
	if (addfprdy = '1') then state := s16080;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16079; end if;
when s16080 => state := s16081; 	--21
	addfpsclr <= '0';
when s16081 => state := s16082; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (786, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16082 => state := s16083; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1510, 12)); -- offset LSB 1462
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s16083 => state := s16084;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1511, 12)); -- offset MSB 1463
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16084 => state := s16085; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16085 => 			--4
	if (fixed2floatrdy = '1') then state := s16086;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16085; end if;
when s16086 => state := s16087; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16087 => 			--6
	if (mulfprdy = '1') then state := s16088;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16087; end if;
when s16088 => state := s16089; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16089 => 			--8
	if (mulfprdy = '1') then state := s16090;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16089; end if;
when s16090 => state := s16091; 	--9
	mulfpsclr <= '0';
when s16091 => state := s16092; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16092 => 			--11
	if (mulfprdy = '1') then state := s16093;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16092; end if;
when s16093 => state := s16094; 	--12
	mulfpsclr <= '0';
when s16094 => state := s16095; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16095 => 			--14
	if (addfprdy = '1') then state := s16096;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16095; end if;
when s16096 => state := s16097; 	--15
	addfpsclr <= '0';
when s16097 => state := s16098; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16098 => 			--17
	if (addfprdy = '1') then state := s16099;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16098; end if;
when s16099 => state := s16100; 	--18
	addfpsclr <= '0';
when s16100 => state := s16101; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16101 => 			--20
	if (addfprdy = '1') then state := s16102;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16101; end if;
when s16102 => state := s16103; 	--21
	addfpsclr <= '0';
when s16103 => state := s16104; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (787, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16104 => state := s16105; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1512, 12)); -- offset LSB 1464
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s16105 => state := s16106;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1513, 12)); -- offset MSB 1465
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16106 => state := s16107; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16107 => 			--4
	if (fixed2floatrdy = '1') then state := s16108;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16107; end if;
when s16108 => state := s16109; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16109 => 			--6
	if (mulfprdy = '1') then state := s16110;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16109; end if;
when s16110 => state := s16111; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16111 => 			--8
	if (mulfprdy = '1') then state := s16112;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16111; end if;
when s16112 => state := s16113; 	--9
	mulfpsclr <= '0';
when s16113 => state := s16114; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16114 => 			--11
	if (mulfprdy = '1') then state := s16115;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16114; end if;
when s16115 => state := s16116; 	--12
	mulfpsclr <= '0';
when s16116 => state := s16117; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16117 => 			--14
	if (addfprdy = '1') then state := s16118;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16117; end if;
when s16118 => state := s16119; 	--15
	addfpsclr <= '0';
when s16119 => state := s16120; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16120 => 			--17
	if (addfprdy = '1') then state := s16121;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16120; end if;
when s16121 => state := s16122; 	--18
	addfpsclr <= '0';
when s16122 => state := s16123; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16123 => 			--20
	if (addfprdy = '1') then state := s16124;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16123; end if;
when s16124 => state := s16125; 	--21
	addfpsclr <= '0';
when s16125 => state := s16126; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (788, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16126 => state := s16127; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1514, 12)); -- offset LSB 1466
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s16127 => state := s16128;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1515, 12)); -- offset MSB 1467
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16128 => state := s16129; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16129 => 			--4
	if (fixed2floatrdy = '1') then state := s16130;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16129; end if;
when s16130 => state := s16131; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16131 => 			--6
	if (mulfprdy = '1') then state := s16132;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16131; end if;
when s16132 => state := s16133; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16133 => 			--8
	if (mulfprdy = '1') then state := s16134;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16133; end if;
when s16134 => state := s16135; 	--9
	mulfpsclr <= '0';
when s16135 => state := s16136; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16136 => 			--11
	if (mulfprdy = '1') then state := s16137;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16136; end if;
when s16137 => state := s16138; 	--12
	mulfpsclr <= '0';
when s16138 => state := s16139; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16139 => 			--14
	if (addfprdy = '1') then state := s16140;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16139; end if;
when s16140 => state := s16141; 	--15
	addfpsclr <= '0';
when s16141 => state := s16142; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16142 => 			--17
	if (addfprdy = '1') then state := s16143;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16142; end if;
when s16143 => state := s16144; 	--18
	addfpsclr <= '0';
when s16144 => state := s16145; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16145 => 			--20
	if (addfprdy = '1') then state := s16146;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16145; end if;
when s16146 => state := s16147; 	--21
	addfpsclr <= '0';
when s16147 => state := s16148; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (789, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16148 => state := s16149; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1516, 12)); -- offset LSB 1468
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s16149 => state := s16150;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1517, 12)); -- offset MSB 1469
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16150 => state := s16151; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16151 => 			--4
	if (fixed2floatrdy = '1') then state := s16152;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16151; end if;
when s16152 => state := s16153; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16153 => 			--6
	if (mulfprdy = '1') then state := s16154;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16153; end if;
when s16154 => state := s16155; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16155 => 			--8
	if (mulfprdy = '1') then state := s16156;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16155; end if;
when s16156 => state := s16157; 	--9
	mulfpsclr <= '0';
when s16157 => state := s16158; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16158 => 			--11
	if (mulfprdy = '1') then state := s16159;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16158; end if;
when s16159 => state := s16160; 	--12
	mulfpsclr <= '0';
when s16160 => state := s16161; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16161 => 			--14
	if (addfprdy = '1') then state := s16162;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16161; end if;
when s16162 => state := s16163; 	--15
	addfpsclr <= '0';
when s16163 => state := s16164; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16164 => 			--17
	if (addfprdy = '1') then state := s16165;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16164; end if;
when s16165 => state := s16166; 	--18
	addfpsclr <= '0';
when s16166 => state := s16167; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16167 => 			--20
	if (addfprdy = '1') then state := s16168;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16167; end if;
when s16168 => state := s16169; 	--21
	addfpsclr <= '0';
when s16169 => state := s16170; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (790, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16170 => state := s16171; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1518, 12)); -- offset LSB 1470
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s16171 => state := s16172;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1519, 12)); -- offset MSB 1471
	addra <= std_logic_vector (to_unsigned (22, 10)); -- OCCrowI 22
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16172 => state := s16173; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16173 => 			--4
	if (fixed2floatrdy = '1') then state := s16174;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16173; end if;
when s16174 => state := s16175; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16175 => 			--6
	if (mulfprdy = '1') then state := s16176;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16175; end if;
when s16176 => state := s16177; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16177 => 			--8
	if (mulfprdy = '1') then state := s16178;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16177; end if;
when s16178 => state := s16179; 	--9
	mulfpsclr <= '0';
when s16179 => state := s16180; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16180 => 			--11
	if (mulfprdy = '1') then state := s16181;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16180; end if;
when s16181 => state := s16182; 	--12
	mulfpsclr <= '0';
when s16182 => state := s16183; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16183 => 			--14
	if (addfprdy = '1') then state := s16184;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16183; end if;
when s16184 => state := s16185; 	--15
	addfpsclr <= '0';
when s16185 => state := s16186; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16186 => 			--17
	if (addfprdy = '1') then state := s16187;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16186; end if;
when s16187 => state := s16188; 	--18
	addfpsclr <= '0';
when s16188 => state := s16189; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16189 => 			--20
	if (addfprdy = '1') then state := s16190;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16189; end if;
when s16190 => state := s16191; 	--21
	addfpsclr <= '0';
when s16191 => state := s16192; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (791, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16192 => state := s16193; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1520, 12)); -- offset LSB 1472
	addra <= std_logic_vector (to_unsigned (24, 10)); -- OCCColumnJ 0
when s16193 => state := s16194;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1521, 12)); -- offset MSB 1473
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16194 => state := s16195; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16195 => 			--4
	if (fixed2floatrdy = '1') then state := s16196;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16195; end if;
when s16196 => state := s16197; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16197 => 			--6
	if (mulfprdy = '1') then state := s16198;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16197; end if;
when s16198 => state := s16199; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16199 => 			--8
	if (mulfprdy = '1') then state := s16200;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16199; end if;
when s16200 => state := s16201; 	--9
	mulfpsclr <= '0';
when s16201 => state := s16202; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16202 => 			--11
	if (mulfprdy = '1') then state := s16203;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16202; end if;
when s16203 => state := s16204; 	--12
	mulfpsclr <= '0';
when s16204 => state := s16205; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16205 => 			--14
	if (addfprdy = '1') then state := s16206;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16205; end if;
when s16206 => state := s16207; 	--15
	addfpsclr <= '0';
when s16207 => state := s16208; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16208 => 			--17
	if (addfprdy = '1') then state := s16209;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16208; end if;
when s16209 => state := s16210; 	--18
	addfpsclr <= '0';
when s16210 => state := s16211; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16211 => 			--20
	if (addfprdy = '1') then state := s16212;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16211; end if;
when s16212 => state := s16213; 	--21
	addfpsclr <= '0';
when s16213 => state := s16214; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (792, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16214 => state := s16215; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1522, 12)); -- offset LSB 1474
	addra <= std_logic_vector (to_unsigned (25, 10)); -- OCCColumnJ 1
when s16215 => state := s16216;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1523, 12)); -- offset MSB 1475
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16216 => state := s16217; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16217 => 			--4
	if (fixed2floatrdy = '1') then state := s16218;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16217; end if;
when s16218 => state := s16219; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16219 => 			--6
	if (mulfprdy = '1') then state := s16220;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16219; end if;
when s16220 => state := s16221; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16221 => 			--8
	if (mulfprdy = '1') then state := s16222;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16221; end if;
when s16222 => state := s16223; 	--9
	mulfpsclr <= '0';
when s16223 => state := s16224; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16224 => 			--11
	if (mulfprdy = '1') then state := s16225;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16224; end if;
when s16225 => state := s16226; 	--12
	mulfpsclr <= '0';
when s16226 => state := s16227; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16227 => 			--14
	if (addfprdy = '1') then state := s16228;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16227; end if;
when s16228 => state := s16229; 	--15
	addfpsclr <= '0';
when s16229 => state := s16230; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16230 => 			--17
	if (addfprdy = '1') then state := s16231;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16230; end if;
when s16231 => state := s16232; 	--18
	addfpsclr <= '0';
when s16232 => state := s16233; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16233 => 			--20
	if (addfprdy = '1') then state := s16234;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16233; end if;
when s16234 => state := s16235; 	--21
	addfpsclr <= '0';
when s16235 => state := s16236; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (793, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16236 => state := s16237; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1524, 12)); -- offset LSB 1476
	addra <= std_logic_vector (to_unsigned (26, 10)); -- OCCColumnJ 2
when s16237 => state := s16238;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1525, 12)); -- offset MSB 1477
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16238 => state := s16239; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16239 => 			--4
	if (fixed2floatrdy = '1') then state := s16240;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16239; end if;
when s16240 => state := s16241; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16241 => 			--6
	if (mulfprdy = '1') then state := s16242;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16241; end if;
when s16242 => state := s16243; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16243 => 			--8
	if (mulfprdy = '1') then state := s16244;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16243; end if;
when s16244 => state := s16245; 	--9
	mulfpsclr <= '0';
when s16245 => state := s16246; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16246 => 			--11
	if (mulfprdy = '1') then state := s16247;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16246; end if;
when s16247 => state := s16248; 	--12
	mulfpsclr <= '0';
when s16248 => state := s16249; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16249 => 			--14
	if (addfprdy = '1') then state := s16250;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16249; end if;
when s16250 => state := s16251; 	--15
	addfpsclr <= '0';
when s16251 => state := s16252; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16252 => 			--17
	if (addfprdy = '1') then state := s16253;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16252; end if;
when s16253 => state := s16254; 	--18
	addfpsclr <= '0';
when s16254 => state := s16255; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16255 => 			--20
	if (addfprdy = '1') then state := s16256;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16255; end if;
when s16256 => state := s16257; 	--21
	addfpsclr <= '0';
when s16257 => state := s16258; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (794, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16258 => state := s16259; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1526, 12)); -- offset LSB 1478
	addra <= std_logic_vector (to_unsigned (27, 10)); -- OCCColumnJ 3
when s16259 => state := s16260;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1527, 12)); -- offset MSB 1479
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16260 => state := s16261; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16261 => 			--4
	if (fixed2floatrdy = '1') then state := s16262;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16261; end if;
when s16262 => state := s16263; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16263 => 			--6
	if (mulfprdy = '1') then state := s16264;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16263; end if;
when s16264 => state := s16265; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16265 => 			--8
	if (mulfprdy = '1') then state := s16266;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16265; end if;
when s16266 => state := s16267; 	--9
	mulfpsclr <= '0';
when s16267 => state := s16268; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16268 => 			--11
	if (mulfprdy = '1') then state := s16269;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16268; end if;
when s16269 => state := s16270; 	--12
	mulfpsclr <= '0';
when s16270 => state := s16271; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16271 => 			--14
	if (addfprdy = '1') then state := s16272;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16271; end if;
when s16272 => state := s16273; 	--15
	addfpsclr <= '0';
when s16273 => state := s16274; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16274 => 			--17
	if (addfprdy = '1') then state := s16275;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16274; end if;
when s16275 => state := s16276; 	--18
	addfpsclr <= '0';
when s16276 => state := s16277; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16277 => 			--20
	if (addfprdy = '1') then state := s16278;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16277; end if;
when s16278 => state := s16279; 	--21
	addfpsclr <= '0';
when s16279 => state := s16280; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (795, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16280 => state := s16281; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1528, 12)); -- offset LSB 1480
	addra <= std_logic_vector (to_unsigned (28, 10)); -- OCCColumnJ 4
when s16281 => state := s16282;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1529, 12)); -- offset MSB 1481
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16282 => state := s16283; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16283 => 			--4
	if (fixed2floatrdy = '1') then state := s16284;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16283; end if;
when s16284 => state := s16285; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16285 => 			--6
	if (mulfprdy = '1') then state := s16286;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16285; end if;
when s16286 => state := s16287; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16287 => 			--8
	if (mulfprdy = '1') then state := s16288;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16287; end if;
when s16288 => state := s16289; 	--9
	mulfpsclr <= '0';
when s16289 => state := s16290; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16290 => 			--11
	if (mulfprdy = '1') then state := s16291;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16290; end if;
when s16291 => state := s16292; 	--12
	mulfpsclr <= '0';
when s16292 => state := s16293; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16293 => 			--14
	if (addfprdy = '1') then state := s16294;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16293; end if;
when s16294 => state := s16295; 	--15
	addfpsclr <= '0';
when s16295 => state := s16296; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16296 => 			--17
	if (addfprdy = '1') then state := s16297;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16296; end if;
when s16297 => state := s16298; 	--18
	addfpsclr <= '0';
when s16298 => state := s16299; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16299 => 			--20
	if (addfprdy = '1') then state := s16300;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16299; end if;
when s16300 => state := s16301; 	--21
	addfpsclr <= '0';
when s16301 => state := s16302; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (796, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16302 => state := s16303; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1530, 12)); -- offset LSB 1482
	addra <= std_logic_vector (to_unsigned (29, 10)); -- OCCColumnJ 5
when s16303 => state := s16304;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1531, 12)); -- offset MSB 1483
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16304 => state := s16305; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16305 => 			--4
	if (fixed2floatrdy = '1') then state := s16306;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16305; end if;
when s16306 => state := s16307; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16307 => 			--6
	if (mulfprdy = '1') then state := s16308;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16307; end if;
when s16308 => state := s16309; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16309 => 			--8
	if (mulfprdy = '1') then state := s16310;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16309; end if;
when s16310 => state := s16311; 	--9
	mulfpsclr <= '0';
when s16311 => state := s16312; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16312 => 			--11
	if (mulfprdy = '1') then state := s16313;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16312; end if;
when s16313 => state := s16314; 	--12
	mulfpsclr <= '0';
when s16314 => state := s16315; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16315 => 			--14
	if (addfprdy = '1') then state := s16316;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16315; end if;
when s16316 => state := s16317; 	--15
	addfpsclr <= '0';
when s16317 => state := s16318; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16318 => 			--17
	if (addfprdy = '1') then state := s16319;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16318; end if;
when s16319 => state := s16320; 	--18
	addfpsclr <= '0';
when s16320 => state := s16321; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16321 => 			--20
	if (addfprdy = '1') then state := s16322;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16321; end if;
when s16322 => state := s16323; 	--21
	addfpsclr <= '0';
when s16323 => state := s16324; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (797, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16324 => state := s16325; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1532, 12)); -- offset LSB 1484
	addra <= std_logic_vector (to_unsigned (30, 10)); -- OCCColumnJ 6
when s16325 => state := s16326;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1533, 12)); -- offset MSB 1485
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16326 => state := s16327; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16327 => 			--4
	if (fixed2floatrdy = '1') then state := s16328;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16327; end if;
when s16328 => state := s16329; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16329 => 			--6
	if (mulfprdy = '1') then state := s16330;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16329; end if;
when s16330 => state := s16331; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16331 => 			--8
	if (mulfprdy = '1') then state := s16332;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16331; end if;
when s16332 => state := s16333; 	--9
	mulfpsclr <= '0';
when s16333 => state := s16334; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16334 => 			--11
	if (mulfprdy = '1') then state := s16335;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16334; end if;
when s16335 => state := s16336; 	--12
	mulfpsclr <= '0';
when s16336 => state := s16337; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16337 => 			--14
	if (addfprdy = '1') then state := s16338;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16337; end if;
when s16338 => state := s16339; 	--15
	addfpsclr <= '0';
when s16339 => state := s16340; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16340 => 			--17
	if (addfprdy = '1') then state := s16341;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16340; end if;
when s16341 => state := s16342; 	--18
	addfpsclr <= '0';
when s16342 => state := s16343; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16343 => 			--20
	if (addfprdy = '1') then state := s16344;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16343; end if;
when s16344 => state := s16345; 	--21
	addfpsclr <= '0';
when s16345 => state := s16346; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (798, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16346 => state := s16347; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1534, 12)); -- offset LSB 1486
	addra <= std_logic_vector (to_unsigned (31, 10)); -- OCCColumnJ 7
when s16347 => state := s16348;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1535, 12)); -- offset MSB 1487
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16348 => state := s16349; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16349 => 			--4
	if (fixed2floatrdy = '1') then state := s16350;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16349; end if;
when s16350 => state := s16351; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16351 => 			--6
	if (mulfprdy = '1') then state := s16352;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16351; end if;
when s16352 => state := s16353; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16353 => 			--8
	if (mulfprdy = '1') then state := s16354;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16353; end if;
when s16354 => state := s16355; 	--9
	mulfpsclr <= '0';
when s16355 => state := s16356; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16356 => 			--11
	if (mulfprdy = '1') then state := s16357;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16356; end if;
when s16357 => state := s16358; 	--12
	mulfpsclr <= '0';
when s16358 => state := s16359; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16359 => 			--14
	if (addfprdy = '1') then state := s16360;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16359; end if;
when s16360 => state := s16361; 	--15
	addfpsclr <= '0';
when s16361 => state := s16362; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16362 => 			--17
	if (addfprdy = '1') then state := s16363;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16362; end if;
when s16363 => state := s16364; 	--18
	addfpsclr <= '0';
when s16364 => state := s16365; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16365 => 			--20
	if (addfprdy = '1') then state := s16366;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16365; end if;
when s16366 => state := s16367; 	--21
	addfpsclr <= '0';
when s16367 => state := s16368; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (799, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16368 => state := s16369; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1536, 12)); -- offset LSB 1488
	addra <= std_logic_vector (to_unsigned (32, 10)); -- OCCColumnJ 8
when s16369 => state := s16370;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1537, 12)); -- offset MSB 1489
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16370 => state := s16371; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16371 => 			--4
	if (fixed2floatrdy = '1') then state := s16372;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16371; end if;
when s16372 => state := s16373; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16373 => 			--6
	if (mulfprdy = '1') then state := s16374;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16373; end if;
when s16374 => state := s16375; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16375 => 			--8
	if (mulfprdy = '1') then state := s16376;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16375; end if;
when s16376 => state := s16377; 	--9
	mulfpsclr <= '0';
when s16377 => state := s16378; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16378 => 			--11
	if (mulfprdy = '1') then state := s16379;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16378; end if;
when s16379 => state := s16380; 	--12
	mulfpsclr <= '0';
when s16380 => state := s16381; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16381 => 			--14
	if (addfprdy = '1') then state := s16382;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16381; end if;
when s16382 => state := s16383; 	--15
	addfpsclr <= '0';
when s16383 => state := s16384; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16384 => 			--17
	if (addfprdy = '1') then state := s16385;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16384; end if;
when s16385 => state := s16386; 	--18
	addfpsclr <= '0';
when s16386 => state := s16387; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16387 => 			--20
	if (addfprdy = '1') then state := s16388;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16387; end if;
when s16388 => state := s16389; 	--21
	addfpsclr <= '0';
when s16389 => state := s16390; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (800, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16390 => state := s16391; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1538, 12)); -- offset LSB 1490
	addra <= std_logic_vector (to_unsigned (33, 10)); -- OCCColumnJ 9
when s16391 => state := s16392;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1539, 12)); -- offset MSB 1491
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16392 => state := s16393; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16393 => 			--4
	if (fixed2floatrdy = '1') then state := s16394;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16393; end if;
when s16394 => state := s16395; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16395 => 			--6
	if (mulfprdy = '1') then state := s16396;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16395; end if;
when s16396 => state := s16397; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16397 => 			--8
	if (mulfprdy = '1') then state := s16398;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16397; end if;
when s16398 => state := s16399; 	--9
	mulfpsclr <= '0';
when s16399 => state := s16400; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16400 => 			--11
	if (mulfprdy = '1') then state := s16401;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16400; end if;
when s16401 => state := s16402; 	--12
	mulfpsclr <= '0';
when s16402 => state := s16403; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16403 => 			--14
	if (addfprdy = '1') then state := s16404;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16403; end if;
when s16404 => state := s16405; 	--15
	addfpsclr <= '0';
when s16405 => state := s16406; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16406 => 			--17
	if (addfprdy = '1') then state := s16407;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16406; end if;
when s16407 => state := s16408; 	--18
	addfpsclr <= '0';
when s16408 => state := s16409; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16409 => 			--20
	if (addfprdy = '1') then state := s16410;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16409; end if;
when s16410 => state := s16411; 	--21
	addfpsclr <= '0';
when s16411 => state := s16412; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (801, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16412 => state := s16413; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1540, 12)); -- offset LSB 1492
	addra <= std_logic_vector (to_unsigned (34, 10)); -- OCCColumnJ 10
when s16413 => state := s16414;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1541, 12)); -- offset MSB 1493
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16414 => state := s16415; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16415 => 			--4
	if (fixed2floatrdy = '1') then state := s16416;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16415; end if;
when s16416 => state := s16417; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16417 => 			--6
	if (mulfprdy = '1') then state := s16418;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16417; end if;
when s16418 => state := s16419; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16419 => 			--8
	if (mulfprdy = '1') then state := s16420;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16419; end if;
when s16420 => state := s16421; 	--9
	mulfpsclr <= '0';
when s16421 => state := s16422; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16422 => 			--11
	if (mulfprdy = '1') then state := s16423;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16422; end if;
when s16423 => state := s16424; 	--12
	mulfpsclr <= '0';
when s16424 => state := s16425; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16425 => 			--14
	if (addfprdy = '1') then state := s16426;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16425; end if;
when s16426 => state := s16427; 	--15
	addfpsclr <= '0';
when s16427 => state := s16428; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16428 => 			--17
	if (addfprdy = '1') then state := s16429;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16428; end if;
when s16429 => state := s16430; 	--18
	addfpsclr <= '0';
when s16430 => state := s16431; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16431 => 			--20
	if (addfprdy = '1') then state := s16432;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16431; end if;
when s16432 => state := s16433; 	--21
	addfpsclr <= '0';
when s16433 => state := s16434; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (802, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16434 => state := s16435; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1542, 12)); -- offset LSB 1494
	addra <= std_logic_vector (to_unsigned (35, 10)); -- OCCColumnJ 11
when s16435 => state := s16436;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1543, 12)); -- offset MSB 1495
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16436 => state := s16437; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16437 => 			--4
	if (fixed2floatrdy = '1') then state := s16438;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16437; end if;
when s16438 => state := s16439; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16439 => 			--6
	if (mulfprdy = '1') then state := s16440;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16439; end if;
when s16440 => state := s16441; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16441 => 			--8
	if (mulfprdy = '1') then state := s16442;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16441; end if;
when s16442 => state := s16443; 	--9
	mulfpsclr <= '0';
when s16443 => state := s16444; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16444 => 			--11
	if (mulfprdy = '1') then state := s16445;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16444; end if;
when s16445 => state := s16446; 	--12
	mulfpsclr <= '0';
when s16446 => state := s16447; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16447 => 			--14
	if (addfprdy = '1') then state := s16448;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16447; end if;
when s16448 => state := s16449; 	--15
	addfpsclr <= '0';
when s16449 => state := s16450; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16450 => 			--17
	if (addfprdy = '1') then state := s16451;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16450; end if;
when s16451 => state := s16452; 	--18
	addfpsclr <= '0';
when s16452 => state := s16453; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16453 => 			--20
	if (addfprdy = '1') then state := s16454;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16453; end if;
when s16454 => state := s16455; 	--21
	addfpsclr <= '0';
when s16455 => state := s16456; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (803, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16456 => state := s16457; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1544, 12)); -- offset LSB 1496
	addra <= std_logic_vector (to_unsigned (36, 10)); -- OCCColumnJ 12
when s16457 => state := s16458;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1545, 12)); -- offset MSB 1497
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16458 => state := s16459; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16459 => 			--4
	if (fixed2floatrdy = '1') then state := s16460;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16459; end if;
when s16460 => state := s16461; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16461 => 			--6
	if (mulfprdy = '1') then state := s16462;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16461; end if;
when s16462 => state := s16463; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16463 => 			--8
	if (mulfprdy = '1') then state := s16464;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16463; end if;
when s16464 => state := s16465; 	--9
	mulfpsclr <= '0';
when s16465 => state := s16466; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16466 => 			--11
	if (mulfprdy = '1') then state := s16467;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16466; end if;
when s16467 => state := s16468; 	--12
	mulfpsclr <= '0';
when s16468 => state := s16469; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16469 => 			--14
	if (addfprdy = '1') then state := s16470;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16469; end if;
when s16470 => state := s16471; 	--15
	addfpsclr <= '0';
when s16471 => state := s16472; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16472 => 			--17
	if (addfprdy = '1') then state := s16473;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16472; end if;
when s16473 => state := s16474; 	--18
	addfpsclr <= '0';
when s16474 => state := s16475; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16475 => 			--20
	if (addfprdy = '1') then state := s16476;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16475; end if;
when s16476 => state := s16477; 	--21
	addfpsclr <= '0';
when s16477 => state := s16478; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (804, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16478 => state := s16479; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1546, 12)); -- offset LSB 1498
	addra <= std_logic_vector (to_unsigned (37, 10)); -- OCCColumnJ 13
when s16479 => state := s16480;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1547, 12)); -- offset MSB 1499
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16480 => state := s16481; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16481 => 			--4
	if (fixed2floatrdy = '1') then state := s16482;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16481; end if;
when s16482 => state := s16483; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16483 => 			--6
	if (mulfprdy = '1') then state := s16484;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16483; end if;
when s16484 => state := s16485; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16485 => 			--8
	if (mulfprdy = '1') then state := s16486;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16485; end if;
when s16486 => state := s16487; 	--9
	mulfpsclr <= '0';
when s16487 => state := s16488; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16488 => 			--11
	if (mulfprdy = '1') then state := s16489;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16488; end if;
when s16489 => state := s16490; 	--12
	mulfpsclr <= '0';
when s16490 => state := s16491; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16491 => 			--14
	if (addfprdy = '1') then state := s16492;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16491; end if;
when s16492 => state := s16493; 	--15
	addfpsclr <= '0';
when s16493 => state := s16494; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16494 => 			--17
	if (addfprdy = '1') then state := s16495;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16494; end if;
when s16495 => state := s16496; 	--18
	addfpsclr <= '0';
when s16496 => state := s16497; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16497 => 			--20
	if (addfprdy = '1') then state := s16498;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16497; end if;
when s16498 => state := s16499; 	--21
	addfpsclr <= '0';
when s16499 => state := s16500; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (805, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16500 => state := s16501; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1548, 12)); -- offset LSB 1500
	addra <= std_logic_vector (to_unsigned (38, 10)); -- OCCColumnJ 14
when s16501 => state := s16502;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1549, 12)); -- offset MSB 1501
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16502 => state := s16503; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16503 => 			--4
	if (fixed2floatrdy = '1') then state := s16504;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16503; end if;
when s16504 => state := s16505; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16505 => 			--6
	if (mulfprdy = '1') then state := s16506;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16505; end if;
when s16506 => state := s16507; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16507 => 			--8
	if (mulfprdy = '1') then state := s16508;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16507; end if;
when s16508 => state := s16509; 	--9
	mulfpsclr <= '0';
when s16509 => state := s16510; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16510 => 			--11
	if (mulfprdy = '1') then state := s16511;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16510; end if;
when s16511 => state := s16512; 	--12
	mulfpsclr <= '0';
when s16512 => state := s16513; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16513 => 			--14
	if (addfprdy = '1') then state := s16514;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16513; end if;
when s16514 => state := s16515; 	--15
	addfpsclr <= '0';
when s16515 => state := s16516; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16516 => 			--17
	if (addfprdy = '1') then state := s16517;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16516; end if;
when s16517 => state := s16518; 	--18
	addfpsclr <= '0';
when s16518 => state := s16519; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16519 => 			--20
	if (addfprdy = '1') then state := s16520;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16519; end if;
when s16520 => state := s16521; 	--21
	addfpsclr <= '0';
when s16521 => state := s16522; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (806, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16522 => state := s16523; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1550, 12)); -- offset LSB 1502
	addra <= std_logic_vector (to_unsigned (39, 10)); -- OCCColumnJ 15
when s16523 => state := s16524;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1551, 12)); -- offset MSB 1503
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16524 => state := s16525; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16525 => 			--4
	if (fixed2floatrdy = '1') then state := s16526;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16525; end if;
when s16526 => state := s16527; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16527 => 			--6
	if (mulfprdy = '1') then state := s16528;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16527; end if;
when s16528 => state := s16529; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16529 => 			--8
	if (mulfprdy = '1') then state := s16530;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16529; end if;
when s16530 => state := s16531; 	--9
	mulfpsclr <= '0';
when s16531 => state := s16532; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16532 => 			--11
	if (mulfprdy = '1') then state := s16533;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16532; end if;
when s16533 => state := s16534; 	--12
	mulfpsclr <= '0';
when s16534 => state := s16535; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16535 => 			--14
	if (addfprdy = '1') then state := s16536;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16535; end if;
when s16536 => state := s16537; 	--15
	addfpsclr <= '0';
when s16537 => state := s16538; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16538 => 			--17
	if (addfprdy = '1') then state := s16539;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16538; end if;
when s16539 => state := s16540; 	--18
	addfpsclr <= '0';
when s16540 => state := s16541; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16541 => 			--20
	if (addfprdy = '1') then state := s16542;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16541; end if;
when s16542 => state := s16543; 	--21
	addfpsclr <= '0';
when s16543 => state := s16544; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (807, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16544 => state := s16545; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1552, 12)); -- offset LSB 1504
	addra <= std_logic_vector (to_unsigned (40, 10)); -- OCCColumnJ 16
when s16545 => state := s16546;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1553, 12)); -- offset MSB 1505
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16546 => state := s16547; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16547 => 			--4
	if (fixed2floatrdy = '1') then state := s16548;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16547; end if;
when s16548 => state := s16549; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16549 => 			--6
	if (mulfprdy = '1') then state := s16550;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16549; end if;
when s16550 => state := s16551; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16551 => 			--8
	if (mulfprdy = '1') then state := s16552;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16551; end if;
when s16552 => state := s16553; 	--9
	mulfpsclr <= '0';
when s16553 => state := s16554; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16554 => 			--11
	if (mulfprdy = '1') then state := s16555;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16554; end if;
when s16555 => state := s16556; 	--12
	mulfpsclr <= '0';
when s16556 => state := s16557; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16557 => 			--14
	if (addfprdy = '1') then state := s16558;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16557; end if;
when s16558 => state := s16559; 	--15
	addfpsclr <= '0';
when s16559 => state := s16560; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16560 => 			--17
	if (addfprdy = '1') then state := s16561;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16560; end if;
when s16561 => state := s16562; 	--18
	addfpsclr <= '0';
when s16562 => state := s16563; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16563 => 			--20
	if (addfprdy = '1') then state := s16564;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16563; end if;
when s16564 => state := s16565; 	--21
	addfpsclr <= '0';
when s16565 => state := s16566; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (808, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16566 => state := s16567; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1554, 12)); -- offset LSB 1506
	addra <= std_logic_vector (to_unsigned (41, 10)); -- OCCColumnJ 17
when s16567 => state := s16568;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1555, 12)); -- offset MSB 1507
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16568 => state := s16569; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16569 => 			--4
	if (fixed2floatrdy = '1') then state := s16570;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16569; end if;
when s16570 => state := s16571; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16571 => 			--6
	if (mulfprdy = '1') then state := s16572;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16571; end if;
when s16572 => state := s16573; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16573 => 			--8
	if (mulfprdy = '1') then state := s16574;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16573; end if;
when s16574 => state := s16575; 	--9
	mulfpsclr <= '0';
when s16575 => state := s16576; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16576 => 			--11
	if (mulfprdy = '1') then state := s16577;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16576; end if;
when s16577 => state := s16578; 	--12
	mulfpsclr <= '0';
when s16578 => state := s16579; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16579 => 			--14
	if (addfprdy = '1') then state := s16580;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16579; end if;
when s16580 => state := s16581; 	--15
	addfpsclr <= '0';
when s16581 => state := s16582; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16582 => 			--17
	if (addfprdy = '1') then state := s16583;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16582; end if;
when s16583 => state := s16584; 	--18
	addfpsclr <= '0';
when s16584 => state := s16585; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16585 => 			--20
	if (addfprdy = '1') then state := s16586;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16585; end if;
when s16586 => state := s16587; 	--21
	addfpsclr <= '0';
when s16587 => state := s16588; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (809, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16588 => state := s16589; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1556, 12)); -- offset LSB 1508
	addra <= std_logic_vector (to_unsigned (42, 10)); -- OCCColumnJ 18
when s16589 => state := s16590;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1557, 12)); -- offset MSB 1509
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16590 => state := s16591; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16591 => 			--4
	if (fixed2floatrdy = '1') then state := s16592;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16591; end if;
when s16592 => state := s16593; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16593 => 			--6
	if (mulfprdy = '1') then state := s16594;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16593; end if;
when s16594 => state := s16595; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16595 => 			--8
	if (mulfprdy = '1') then state := s16596;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16595; end if;
when s16596 => state := s16597; 	--9
	mulfpsclr <= '0';
when s16597 => state := s16598; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16598 => 			--11
	if (mulfprdy = '1') then state := s16599;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16598; end if;
when s16599 => state := s16600; 	--12
	mulfpsclr <= '0';
when s16600 => state := s16601; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16601 => 			--14
	if (addfprdy = '1') then state := s16602;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16601; end if;
when s16602 => state := s16603; 	--15
	addfpsclr <= '0';
when s16603 => state := s16604; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16604 => 			--17
	if (addfprdy = '1') then state := s16605;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16604; end if;
when s16605 => state := s16606; 	--18
	addfpsclr <= '0';
when s16606 => state := s16607; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16607 => 			--20
	if (addfprdy = '1') then state := s16608;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16607; end if;
when s16608 => state := s16609; 	--21
	addfpsclr <= '0';
when s16609 => state := s16610; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (810, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16610 => state := s16611; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1558, 12)); -- offset LSB 1510
	addra <= std_logic_vector (to_unsigned (43, 10)); -- OCCColumnJ 19
when s16611 => state := s16612;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1559, 12)); -- offset MSB 1511
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16612 => state := s16613; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16613 => 			--4
	if (fixed2floatrdy = '1') then state := s16614;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16613; end if;
when s16614 => state := s16615; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16615 => 			--6
	if (mulfprdy = '1') then state := s16616;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16615; end if;
when s16616 => state := s16617; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16617 => 			--8
	if (mulfprdy = '1') then state := s16618;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16617; end if;
when s16618 => state := s16619; 	--9
	mulfpsclr <= '0';
when s16619 => state := s16620; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16620 => 			--11
	if (mulfprdy = '1') then state := s16621;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16620; end if;
when s16621 => state := s16622; 	--12
	mulfpsclr <= '0';
when s16622 => state := s16623; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16623 => 			--14
	if (addfprdy = '1') then state := s16624;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16623; end if;
when s16624 => state := s16625; 	--15
	addfpsclr <= '0';
when s16625 => state := s16626; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16626 => 			--17
	if (addfprdy = '1') then state := s16627;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16626; end if;
when s16627 => state := s16628; 	--18
	addfpsclr <= '0';
when s16628 => state := s16629; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16629 => 			--20
	if (addfprdy = '1') then state := s16630;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16629; end if;
when s16630 => state := s16631; 	--21
	addfpsclr <= '0';
when s16631 => state := s16632; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (811, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16632 => state := s16633; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1560, 12)); -- offset LSB 1512
	addra <= std_logic_vector (to_unsigned (44, 10)); -- OCCColumnJ 20
when s16633 => state := s16634;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1561, 12)); -- offset MSB 1513
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16634 => state := s16635; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16635 => 			--4
	if (fixed2floatrdy = '1') then state := s16636;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16635; end if;
when s16636 => state := s16637; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16637 => 			--6
	if (mulfprdy = '1') then state := s16638;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16637; end if;
when s16638 => state := s16639; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16639 => 			--8
	if (mulfprdy = '1') then state := s16640;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16639; end if;
when s16640 => state := s16641; 	--9
	mulfpsclr <= '0';
when s16641 => state := s16642; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16642 => 			--11
	if (mulfprdy = '1') then state := s16643;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16642; end if;
when s16643 => state := s16644; 	--12
	mulfpsclr <= '0';
when s16644 => state := s16645; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16645 => 			--14
	if (addfprdy = '1') then state := s16646;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16645; end if;
when s16646 => state := s16647; 	--15
	addfpsclr <= '0';
when s16647 => state := s16648; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16648 => 			--17
	if (addfprdy = '1') then state := s16649;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16648; end if;
when s16649 => state := s16650; 	--18
	addfpsclr <= '0';
when s16650 => state := s16651; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16651 => 			--20
	if (addfprdy = '1') then state := s16652;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16651; end if;
when s16652 => state := s16653; 	--21
	addfpsclr <= '0';
when s16653 => state := s16654; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (812, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16654 => state := s16655; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1562, 12)); -- offset LSB 1514
	addra <= std_logic_vector (to_unsigned (45, 10)); -- OCCColumnJ 21
when s16655 => state := s16656;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1563, 12)); -- offset MSB 1515
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16656 => state := s16657; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16657 => 			--4
	if (fixed2floatrdy = '1') then state := s16658;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16657; end if;
when s16658 => state := s16659; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16659 => 			--6
	if (mulfprdy = '1') then state := s16660;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16659; end if;
when s16660 => state := s16661; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16661 => 			--8
	if (mulfprdy = '1') then state := s16662;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16661; end if;
when s16662 => state := s16663; 	--9
	mulfpsclr <= '0';
when s16663 => state := s16664; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16664 => 			--11
	if (mulfprdy = '1') then state := s16665;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16664; end if;
when s16665 => state := s16666; 	--12
	mulfpsclr <= '0';
when s16666 => state := s16667; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16667 => 			--14
	if (addfprdy = '1') then state := s16668;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16667; end if;
when s16668 => state := s16669; 	--15
	addfpsclr <= '0';
when s16669 => state := s16670; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16670 => 			--17
	if (addfprdy = '1') then state := s16671;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16670; end if;
when s16671 => state := s16672; 	--18
	addfpsclr <= '0';
when s16672 => state := s16673; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16673 => 			--20
	if (addfprdy = '1') then state := s16674;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16673; end if;
when s16674 => state := s16675; 	--21
	addfpsclr <= '0';
when s16675 => state := s16676; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (813, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16676 => state := s16677; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1564, 12)); -- offset LSB 1516
	addra <= std_logic_vector (to_unsigned (46, 10)); -- OCCColumnJ 22
when s16677 => state := s16678;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1565, 12)); -- offset MSB 1517
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16678 => state := s16679; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16679 => 			--4
	if (fixed2floatrdy = '1') then state := s16680;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16679; end if;
when s16680 => state := s16681; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16681 => 			--6
	if (mulfprdy = '1') then state := s16682;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16681; end if;
when s16682 => state := s16683; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16683 => 			--8
	if (mulfprdy = '1') then state := s16684;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16683; end if;
when s16684 => state := s16685; 	--9
	mulfpsclr <= '0';
when s16685 => state := s16686; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16686 => 			--11
	if (mulfprdy = '1') then state := s16687;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16686; end if;
when s16687 => state := s16688; 	--12
	mulfpsclr <= '0';
when s16688 => state := s16689; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16689 => 			--14
	if (addfprdy = '1') then state := s16690;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16689; end if;
when s16690 => state := s16691; 	--15
	addfpsclr <= '0';
when s16691 => state := s16692; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16692 => 			--17
	if (addfprdy = '1') then state := s16693;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16692; end if;
when s16693 => state := s16694; 	--18
	addfpsclr <= '0';
when s16694 => state := s16695; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16695 => 			--20
	if (addfprdy = '1') then state := s16696;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16695; end if;
when s16696 => state := s16697; 	--21
	addfpsclr <= '0';
when s16697 => state := s16698; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (814, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16698 => state := s16699; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1566, 12)); -- offset LSB 1518
	addra <= std_logic_vector (to_unsigned (47, 10)); -- OCCColumnJ 23
when s16699 => state := s16700;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1567, 12)); -- offset MSB 1519
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16700 => state := s16701; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16701 => 			--4
	if (fixed2floatrdy = '1') then state := s16702;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16701; end if;
when s16702 => state := s16703; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16703 => 			--6
	if (mulfprdy = '1') then state := s16704;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16703; end if;
when s16704 => state := s16705; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16705 => 			--8
	if (mulfprdy = '1') then state := s16706;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16705; end if;
when s16706 => state := s16707; 	--9
	mulfpsclr <= '0';
when s16707 => state := s16708; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16708 => 			--11
	if (mulfprdy = '1') then state := s16709;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16708; end if;
when s16709 => state := s16710; 	--12
	mulfpsclr <= '0';
when s16710 => state := s16711; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16711 => 			--14
	if (addfprdy = '1') then state := s16712;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16711; end if;
when s16712 => state := s16713; 	--15
	addfpsclr <= '0';
when s16713 => state := s16714; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16714 => 			--17
	if (addfprdy = '1') then state := s16715;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16714; end if;
when s16715 => state := s16716; 	--18
	addfpsclr <= '0';
when s16716 => state := s16717; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16717 => 			--20
	if (addfprdy = '1') then state := s16718;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16717; end if;
when s16718 => state := s16719; 	--21
	addfpsclr <= '0';
when s16719 => state := s16720; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (815, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16720 => state := s16721; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1568, 12)); -- offset LSB 1520
	addra <= std_logic_vector (to_unsigned (48, 10)); -- OCCColumnJ 24
when s16721 => state := s16722;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1569, 12)); -- offset MSB 1521
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16722 => state := s16723; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16723 => 			--4
	if (fixed2floatrdy = '1') then state := s16724;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16723; end if;
when s16724 => state := s16725; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16725 => 			--6
	if (mulfprdy = '1') then state := s16726;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16725; end if;
when s16726 => state := s16727; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16727 => 			--8
	if (mulfprdy = '1') then state := s16728;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16727; end if;
when s16728 => state := s16729; 	--9
	mulfpsclr <= '0';
when s16729 => state := s16730; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16730 => 			--11
	if (mulfprdy = '1') then state := s16731;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16730; end if;
when s16731 => state := s16732; 	--12
	mulfpsclr <= '0';
when s16732 => state := s16733; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16733 => 			--14
	if (addfprdy = '1') then state := s16734;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16733; end if;
when s16734 => state := s16735; 	--15
	addfpsclr <= '0';
when s16735 => state := s16736; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16736 => 			--17
	if (addfprdy = '1') then state := s16737;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16736; end if;
when s16737 => state := s16738; 	--18
	addfpsclr <= '0';
when s16738 => state := s16739; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16739 => 			--20
	if (addfprdy = '1') then state := s16740;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16739; end if;
when s16740 => state := s16741; 	--21
	addfpsclr <= '0';
when s16741 => state := s16742; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (816, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16742 => state := s16743; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1570, 12)); -- offset LSB 1522
	addra <= std_logic_vector (to_unsigned (49, 10)); -- OCCColumnJ 25
when s16743 => state := s16744;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1571, 12)); -- offset MSB 1523
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16744 => state := s16745; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16745 => 			--4
	if (fixed2floatrdy = '1') then state := s16746;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16745; end if;
when s16746 => state := s16747; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16747 => 			--6
	if (mulfprdy = '1') then state := s16748;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16747; end if;
when s16748 => state := s16749; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16749 => 			--8
	if (mulfprdy = '1') then state := s16750;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16749; end if;
when s16750 => state := s16751; 	--9
	mulfpsclr <= '0';
when s16751 => state := s16752; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16752 => 			--11
	if (mulfprdy = '1') then state := s16753;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16752; end if;
when s16753 => state := s16754; 	--12
	mulfpsclr <= '0';
when s16754 => state := s16755; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16755 => 			--14
	if (addfprdy = '1') then state := s16756;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16755; end if;
when s16756 => state := s16757; 	--15
	addfpsclr <= '0';
when s16757 => state := s16758; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16758 => 			--17
	if (addfprdy = '1') then state := s16759;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16758; end if;
when s16759 => state := s16760; 	--18
	addfpsclr <= '0';
when s16760 => state := s16761; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16761 => 			--20
	if (addfprdy = '1') then state := s16762;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16761; end if;
when s16762 => state := s16763; 	--21
	addfpsclr <= '0';
when s16763 => state := s16764; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (817, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16764 => state := s16765; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1572, 12)); -- offset LSB 1524
	addra <= std_logic_vector (to_unsigned (50, 10)); -- OCCColumnJ 26
when s16765 => state := s16766;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1573, 12)); -- offset MSB 1525
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16766 => state := s16767; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16767 => 			--4
	if (fixed2floatrdy = '1') then state := s16768;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16767; end if;
when s16768 => state := s16769; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16769 => 			--6
	if (mulfprdy = '1') then state := s16770;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16769; end if;
when s16770 => state := s16771; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16771 => 			--8
	if (mulfprdy = '1') then state := s16772;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16771; end if;
when s16772 => state := s16773; 	--9
	mulfpsclr <= '0';
when s16773 => state := s16774; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16774 => 			--11
	if (mulfprdy = '1') then state := s16775;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16774; end if;
when s16775 => state := s16776; 	--12
	mulfpsclr <= '0';
when s16776 => state := s16777; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16777 => 			--14
	if (addfprdy = '1') then state := s16778;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16777; end if;
when s16778 => state := s16779; 	--15
	addfpsclr <= '0';
when s16779 => state := s16780; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16780 => 			--17
	if (addfprdy = '1') then state := s16781;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16780; end if;
when s16781 => state := s16782; 	--18
	addfpsclr <= '0';
when s16782 => state := s16783; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16783 => 			--20
	if (addfprdy = '1') then state := s16784;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16783; end if;
when s16784 => state := s16785; 	--21
	addfpsclr <= '0';
when s16785 => state := s16786; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (818, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16786 => state := s16787; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1574, 12)); -- offset LSB 1526
	addra <= std_logic_vector (to_unsigned (51, 10)); -- OCCColumnJ 27
when s16787 => state := s16788;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1575, 12)); -- offset MSB 1527
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16788 => state := s16789; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16789 => 			--4
	if (fixed2floatrdy = '1') then state := s16790;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16789; end if;
when s16790 => state := s16791; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16791 => 			--6
	if (mulfprdy = '1') then state := s16792;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16791; end if;
when s16792 => state := s16793; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16793 => 			--8
	if (mulfprdy = '1') then state := s16794;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16793; end if;
when s16794 => state := s16795; 	--9
	mulfpsclr <= '0';
when s16795 => state := s16796; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16796 => 			--11
	if (mulfprdy = '1') then state := s16797;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16796; end if;
when s16797 => state := s16798; 	--12
	mulfpsclr <= '0';
when s16798 => state := s16799; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16799 => 			--14
	if (addfprdy = '1') then state := s16800;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16799; end if;
when s16800 => state := s16801; 	--15
	addfpsclr <= '0';
when s16801 => state := s16802; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16802 => 			--17
	if (addfprdy = '1') then state := s16803;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16802; end if;
when s16803 => state := s16804; 	--18
	addfpsclr <= '0';
when s16804 => state := s16805; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16805 => 			--20
	if (addfprdy = '1') then state := s16806;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16805; end if;
when s16806 => state := s16807; 	--21
	addfpsclr <= '0';
when s16807 => state := s16808; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (819, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16808 => state := s16809; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1576, 12)); -- offset LSB 1528
	addra <= std_logic_vector (to_unsigned (52, 10)); -- OCCColumnJ 28
when s16809 => state := s16810;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1577, 12)); -- offset MSB 1529
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16810 => state := s16811; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16811 => 			--4
	if (fixed2floatrdy = '1') then state := s16812;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16811; end if;
when s16812 => state := s16813; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16813 => 			--6
	if (mulfprdy = '1') then state := s16814;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16813; end if;
when s16814 => state := s16815; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16815 => 			--8
	if (mulfprdy = '1') then state := s16816;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16815; end if;
when s16816 => state := s16817; 	--9
	mulfpsclr <= '0';
when s16817 => state := s16818; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16818 => 			--11
	if (mulfprdy = '1') then state := s16819;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16818; end if;
when s16819 => state := s16820; 	--12
	mulfpsclr <= '0';
when s16820 => state := s16821; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16821 => 			--14
	if (addfprdy = '1') then state := s16822;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16821; end if;
when s16822 => state := s16823; 	--15
	addfpsclr <= '0';
when s16823 => state := s16824; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16824 => 			--17
	if (addfprdy = '1') then state := s16825;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16824; end if;
when s16825 => state := s16826; 	--18
	addfpsclr <= '0';
when s16826 => state := s16827; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16827 => 			--20
	if (addfprdy = '1') then state := s16828;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16827; end if;
when s16828 => state := s16829; 	--21
	addfpsclr <= '0';
when s16829 => state := s16830; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (820, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16830 => state := s16831; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1578, 12)); -- offset LSB 1530
	addra <= std_logic_vector (to_unsigned (53, 10)); -- OCCColumnJ 29
when s16831 => state := s16832;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1579, 12)); -- offset MSB 1531
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16832 => state := s16833; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16833 => 			--4
	if (fixed2floatrdy = '1') then state := s16834;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16833; end if;
when s16834 => state := s16835; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16835 => 			--6
	if (mulfprdy = '1') then state := s16836;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16835; end if;
when s16836 => state := s16837; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16837 => 			--8
	if (mulfprdy = '1') then state := s16838;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16837; end if;
when s16838 => state := s16839; 	--9
	mulfpsclr <= '0';
when s16839 => state := s16840; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16840 => 			--11
	if (mulfprdy = '1') then state := s16841;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16840; end if;
when s16841 => state := s16842; 	--12
	mulfpsclr <= '0';
when s16842 => state := s16843; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16843 => 			--14
	if (addfprdy = '1') then state := s16844;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16843; end if;
when s16844 => state := s16845; 	--15
	addfpsclr <= '0';
when s16845 => state := s16846; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16846 => 			--17
	if (addfprdy = '1') then state := s16847;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16846; end if;
when s16847 => state := s16848; 	--18
	addfpsclr <= '0';
when s16848 => state := s16849; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16849 => 			--20
	if (addfprdy = '1') then state := s16850;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16849; end if;
when s16850 => state := s16851; 	--21
	addfpsclr <= '0';
when s16851 => state := s16852; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (821, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16852 => state := s16853; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1580, 12)); -- offset LSB 1532
	addra <= std_logic_vector (to_unsigned (54, 10)); -- OCCColumnJ 30
when s16853 => state := s16854;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1581, 12)); -- offset MSB 1533
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16854 => state := s16855; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16855 => 			--4
	if (fixed2floatrdy = '1') then state := s16856;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16855; end if;
when s16856 => state := s16857; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16857 => 			--6
	if (mulfprdy = '1') then state := s16858;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16857; end if;
when s16858 => state := s16859; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16859 => 			--8
	if (mulfprdy = '1') then state := s16860;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16859; end if;
when s16860 => state := s16861; 	--9
	mulfpsclr <= '0';
when s16861 => state := s16862; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16862 => 			--11
	if (mulfprdy = '1') then state := s16863;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16862; end if;
when s16863 => state := s16864; 	--12
	mulfpsclr <= '0';
when s16864 => state := s16865; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16865 => 			--14
	if (addfprdy = '1') then state := s16866;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16865; end if;
when s16866 => state := s16867; 	--15
	addfpsclr <= '0';
when s16867 => state := s16868; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16868 => 			--17
	if (addfprdy = '1') then state := s16869;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16868; end if;
when s16869 => state := s16870; 	--18
	addfpsclr <= '0';
when s16870 => state := s16871; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16871 => 			--20
	if (addfprdy = '1') then state := s16872;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16871; end if;
when s16872 => state := s16873; 	--21
	addfpsclr <= '0';
when s16873 => state := s16874; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (822, 10)); -- vOffset_ft
	dia <= vOffset_ft;

when s16874 => state := s16875; 	--1
	write_enable <= '0';
	i2c_mem_addra <= std_logic_vector (to_unsigned (1582, 12)); -- offset LSB 1534
	addra <= std_logic_vector (to_unsigned (55, 10)); -- OCCColumnJ 31
when s16875 => state := s16876;	--2
	i2c_mem_addra <= std_logic_vector (to_unsigned (1583, 12)); -- offset MSB 1535
	addra <= std_logic_vector (to_unsigned (23, 10)); -- OCCrowI 23
	vOCCColumnJ := doa;
	vOffset (7 downto 0) := i2c_mem_douta;
when s16876 => state := s16877; 	--3
	vOCCRowI := doa;
	vOffset (15 downto 8) := i2c_mem_douta;
	vOffset_sf := resize (to_sfixed (vOffset, eeprom16sf), vOffset_sf);
	fixed2floatce <= '1';
	fixed2floatond <= '1';
	fixed2floata <= 
	to_slv (to_sfixed (to_slv (vOffset_sf (fracas'high downto fracas'low)), fracas))&
	to_slv (to_sfixed (to_slv (vOffset_sf (fracbs'high downto fracbs'low)), fracbs));
when s16877 => 			--4
	if (fixed2floatrdy = '1') then state := s16878;
		vOffset_ft := fixed2floatr;
		fixed2floatce <= '0';
		fixed2floatond <= '0';
		fixed2floatsclr <= '1';
	else state := s16877; end if;
when s16878 => state := s16879; 	--5
	fixed2floatsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOffset_ft;
	mulfpb <= voccRemScale;
	mulfpond <= '1';
when s16879 => 			--6
	if (mulfprdy = '1') then state := s16880;
		vOffset_ft := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16879; end if;
when s16880 => state := s16881; 	--7
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCColumnJ;
	mulfpb <= voccColumnScale;
	mulfpond <= '1';
when s16881 => 			--8
	if (mulfprdy = '1') then state := s16882;
		vOCCColumnJ := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16881; end if;
when s16882 => state := s16883; 	--9
	mulfpsclr <= '0';
when s16883 => state := s16884; 	--10
	mulfpsclr <= '0';
	mulfpce <= '1';
	mulfpa <= vOCCRowI;
	mulfpb <= voccRowScale;
	mulfpond <= '1';
when s16884 => 			--11
	if (mulfprdy = '1') then state := s16885;
		vOCCRowI := mulfpr;
		mulfpce <= '0';
		mulfpond <= '0';
		mulfpsclr <= '1';
	else state := s16884; end if;
when s16885 => state := s16886; 	--12
	mulfpsclr <= '0';
when s16886 => state := s16887; 	--13
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCColumnJ;
	addfpond <= '1';
when s16887 => 			--14
	if (addfprdy = '1') then state := s16888;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16887; end if;
when s16888 => state := s16889; 	--15
	addfpsclr <= '0';
when s16889 => state := s16890; 	--16
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOCCRowI;
	addfpond <= '1';
when s16890 => 			--17
	if (addfprdy = '1') then state := s16891;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16890; end if;
when s16891 => state := s16892; 	--18
	addfpsclr <= '0';
when s16892 => state := s16893; 	--19
	addfpsclr <= '0';
	addfpce <= '1';
	addfpa <= vOffset_ft;
	addfpb <= vOffsetAverage;
	addfpond <= '1';
when s16893 => 			--20
	if (addfprdy = '1') then state := s16894;
		vOffset_ft := addfpr;
		addfpce <= '0';
		addfpond <= '0';
		addfpsclr <= '1';
	else state := s16893; end if;
when s16894 => state := s16895; 	--21
	addfpsclr <= '0';
when s16895 => state := ending; 	--22
	write_enable <= '1';
	addra <= std_logic_vector (to_unsigned (823, 10)); -- vOffset_ft
	dia <= vOffset_ft;


				when ending => state := idle;
					rdy <= '1';
				when others => null;
			end case;
--			stemp1 <= temp1;
		end if;
	end if;
end process p0;

inst_mem_occ : mem_ramb16_s36_x2
GENERIC MAP (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000" -- start 0's
)
PORT MAP (
DO => doa,
DOP => open,
ADDR => mux_addr,
CLK => i_clock,
DI => mux_dia,
DIP => (others => '0'),
EN => '1',
SSR => i_reset,
WE => write_enable
);

mulfpclk <= i_clock;
inst_mulfp_acc : mulfp
PORT MAP (
a => mulfpa,
b => mulfpb,
operation_nd => mulfpond,
clk => mulfpclk,
sclr => mulfpsclr,
ce => mulfpce,
result => mulfpr,
rdy => mulfprdy
);

addfpclk <= i_clock;
inst_addfp_acc : addfp
PORT MAP (
a => addfpa,
b => addfpb,
operation_nd => addfpond,
clk => addfpclk,
sclr => addfpsclr,
ce => addfpce,
result => addfpr,
rdy => addfprdy
);

--INIT_7f => X"41700000 41600000 41500000 41400000 41300000 41200000 41100000 41000000", -- unsigned 0-15 for accremscale,accrowscale,acccolscale
--INIT_7e => X"40e00000 40c00000 40a00000 40800000 40400000 40000000 3f800000 22000000",
with nibble1 select out_nibble1 <= -- x - occremscale,occrowscale,occcolscale
x"00000000" when x"0", x"3f800000" when x"1", x"40000000" when x"2", x"40400000" when x"3",
x"40800000" when x"4", x"40a00000" when x"5", x"40c00000" when x"6", x"40e00000" when x"7",
x"41000000" when x"8", x"41100000" when x"9", x"41200000" when x"a", x"41300000" when x"b",
x"41400000" when x"c", x"41500000" when x"d", x"41600000" when x"e", x"41700000" when x"f",
x"00000000" when others;

with nibble2 select out_nibble2 <= -- >7,-16 - rows1-24,cols1-32
x"00000000" when x"0", x"3f800000" when x"1", x"40000000" when x"2", x"40400000" when x"3",
x"40800000" when x"4", x"40a00000" when x"5", x"40c00000" when x"6", x"40e00000" when x"7",
x"c1000000" when x"8", x"c0e00000" when x"9", x"c0c00000" when x"a", x"c0a00000" when x"b",
x"c0800000" when x"c", x"c0400000" when x"d", x"c0000000" when x"e", x"bf800000" when x"f",
x"00000000" when others;

with nibble3 select out_nibble3 <= -- >31,-64 - offset raw
x"40e00000" when "000111",x"40c00000" when "000110",x"40a00000" when "000101",x"40800000" when "000100",x"40400000" when "000011",x"40000000" when "000010",x"3f800000" when "000001",x"22000000" when "000000",
x"41700000" when "001111",x"41600000" when "001110",x"41500000" when "001101",x"41400000" when "001100",x"41300000" when "001011",x"41200000" when "001010",x"41100000" when "001001",x"41000000" when "001000",
x"41b80000" when "010111",x"41b00000" when "010110",x"41a80000" when "010101",x"41a00000" when "010100",x"41980000" when "010011",x"41900000" when "010010",x"41880000" when "010001",x"41800000" when "010000",
x"41f80000" when "011111",x"41f00000" when "011110",x"41e80000" when "011101",x"41e00000" when "011100",x"41d80000" when "011011",x"41d00000" when "011010",x"41c80000" when "011001",x"41c00000" when "011000",
x"c1c80000" when "100111",x"c1d00000" when "100110",x"c1d80000" when "100101",x"c1e00000" when "100100",x"c1e80000" when "100011",x"c1f00000" when "100010",x"c1f80000" when "100001",x"c2000000" when "100000",
x"c1880000" when "101111",x"c1900000" when "101110",x"c1980000" when "101101",x"c1a00000" when "101100",x"c1a80000" when "101011",x"c1b00000" when "101010",x"c1b80000" when "101001",x"c1c00000" when "101000",
x"c1100000" when "110111",x"c1200000" when "110110",x"c1300000" when "110101",x"c1400000" when "110100",x"c1500000" when "110011",x"c1600000" when "110010",x"c1700000" when "110001",x"c1800000" when "110000",
x"bf800000" when "111111",x"c0000000" when "111110",x"c0400000" when "111101",x"c0800000" when "111100",x"c0a00000" when "111011",x"c0c00000" when "111010",x"c0e00000" when "111001",x"c1000000" when "111000",
x"22000000" when others;

--INIT_01 => X"47000000 46800000 46000000 45800000 45000000 44800000 44000000 43800000",
--INIT_00 => X"43000000 42800000 42000000 41800000 41000000 40800000 40000000 3f800000",
with nibble4 select out_nibble4 <= -- 2^x unsigned 0-15
x"3f800000" when x"0", x"40000000" when x"1", x"40800000" when x"2", x"41000000" when x"3",
x"41800000" when x"4", x"42000000" when x"5", x"42800000" when x"6", x"43000000" when x"7",
x"43800000" when x"8", x"44000000" when x"9", x"44800000" when x"a", x"45000000" when x"b",
x"45800000" when x"c", x"46000000" when x"d", x"46800000" when x"e", x"47000000" when x"f",
x"00000000" when others;

fixed2floatclk <= i_clock;
inst_ff2 : fixed2float
PORT MAP (
a => fixed2floata,
operation_nd => fixed2floatond,
clk => fixed2floatclk,
sclr => fixed2floatsclr,
ce => fixed2floatce,
result => fixed2floatr,
rdy => fixed2floatrdy
);

end Behavioral;

