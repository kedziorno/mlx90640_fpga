library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.p_package1_constants.all;

package p_package1 is


end p_package1;

package body p_package1 is

 
end p_package1;
