----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:08:52 02/06/2023 
-- Design Name: 
-- Module Name:    mem_signed1024 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mem_signed1024 is
port (
i_clock : in std_logic;
i_reset : in std_logic;
i_value : in std_logic_vector (9 downto 0); -- input hex from 0 to 1024
o_value : out std_logic_vector (31 downto 0) -- output signed -512 to 511 in SP float
);
end mem_signed1024;

architecture Behavioral of mem_signed1024 is

COMPONENT mem_ramb16_s36_x2
generic (
INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0a : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0b : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0c : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0d : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0e : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
INITP_0f : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
);
PORT(
DO : OUT  std_logic_vector(31 downto 0);
DOP : OUT  std_logic_vector(3 downto 0);
ADDR : IN  std_logic_vector(9 downto 0);
CLK : IN  std_logic;
DI : IN  std_logic_vector(31 downto 0);
DIP : IN  std_logic_vector(3 downto 0);
EN : IN  std_logic;
SSR : IN  std_logic;
WE : IN  std_logic
);
END COMPONENT mem_ramb16_s36_x2;

begin

inst_signed1024 : mem_ramb16_s36_x2 
GENERIC MAP (
INIT_00 => X"40e0000040c0000040a000004080000040400000400000003f80000000000000",       
INIT_01 => X"4170000041600000415000004140000041300000412000004110000041000000",
INIT_02 => X"41b8000041b0000041a8000041a0000041980000419000004188000041800000",
INIT_03 => X"41f8000041f0000041e8000041e0000041d8000041d0000041c8000041c00000",
INIT_04 => X"421c0000421800004214000042100000420c0000420800004204000042000000",
INIT_05 => X"423c0000423800004234000042300000422c0000422800004224000042200000",
INIT_06 => X"425c0000425800004254000042500000424c0000424800004244000042400000",
INIT_07 => X"427c0000427800004274000042700000426c0000426800004264000042600000",
INIT_08 => X"428e0000428c0000428a00004288000042860000428400004282000042800000",
INIT_09 => X"429e0000429c0000429a00004298000042960000429400004292000042900000",
INIT_0a => X"42ae000042ac000042aa000042a8000042a6000042a4000042a2000042a00000",
INIT_0b => X"42be000042bc000042ba000042b8000042b6000042b4000042b2000042b00000",
INIT_0c => X"42ce000042cc000042ca000042c8000042c6000042c4000042c2000042c00000",
INIT_0d => X"42de000042dc000042da000042d8000042d6000042d4000042d2000042d00000",
INIT_0e => X"42ee000042ec000042ea000042e8000042e6000042e4000042e2000042e00000",
INIT_0f => X"42fe000042fc000042fa000042f8000042f6000042f4000042f2000042f00000",
INIT_10 => X"4307000043060000430500004304000043030000430200004301000043000000",
INIT_11 => X"430f0000430e0000430d0000430c0000430b0000430a00004309000043080000",
INIT_12 => X"4317000043160000431500004314000043130000431200004311000043100000",
INIT_13 => X"431f0000431e0000431d0000431c0000431b0000431a00004319000043180000",
INIT_14 => X"4327000043260000432500004324000043230000432200004321000043200000",
INIT_15 => X"432f0000432e0000432d0000432c0000432b0000432a00004329000043280000",
INIT_16 => X"4337000043360000433500004334000043330000433200004331000043300000",
INIT_17 => X"433f0000433e0000433d0000433c0000433b0000433a00004339000043380000",
INIT_18 => X"4347000043460000434500004344000043430000434200004341000043400000",
INIT_19 => X"434f0000434e0000434d0000434c0000434b0000434a00004349000043480000",
INIT_1a => X"4357000043560000435500004354000043530000435200004351000043500000",
INIT_1b => X"435f0000435e0000435d0000435c0000435b0000435a00004359000043580000",
INIT_1c => X"4367000043660000436500004364000043630000436200004361000043600000",
INIT_1d => X"436f0000436e0000436d0000436c0000436b0000436a00004369000043680000",
INIT_1e => X"4377000043760000437500004374000043730000437200004371000043700000",
INIT_1f => X"437f0000437e0000437d0000437c0000437b0000437a00004379000043780000",
INIT_20 => X"4383800043830000438280004382000043818000438100004380800043800000",
INIT_21 => X"4387800043870000438680004386000043858000438500004384800043840000",
INIT_22 => X"438b8000438b0000438a8000438a000043898000438900004388800043880000",
INIT_23 => X"438f8000438f0000438e8000438e0000438d8000438d0000438c8000438c0000",
INIT_24 => X"4393800043930000439280004392000043918000439100004390800043900000",
INIT_25 => X"4397800043970000439680004396000043958000439500004394800043940000",
INIT_26 => X"439b8000439b0000439a8000439a000043998000439900004398800043980000",
INIT_27 => X"439f8000439f0000439e8000439e0000439d8000439d0000439c8000439c0000",
INIT_28 => X"43a3800043a3000043a2800043a2000043a1800043a1000043a0800043a00000",
INIT_29 => X"43a7800043a7000043a6800043a6000043a5800043a5000043a4800043a40000",
INIT_2a => X"43ab800043ab000043aa800043aa000043a9800043a9000043a8800043a80000",
INIT_2b => X"43af800043af000043ae800043ae000043ad800043ad000043ac800043ac0000",
INIT_2c => X"43b3800043b3000043b2800043b2000043b1800043b1000043b0800043b00000",
INIT_2d => X"43b7800043b7000043b6800043b6000043b5800043b5000043b4800043b40000",
INIT_2e => X"43bb800043bb000043ba800043ba000043b9800043b9000043b8800043b80000",
INIT_2f => X"43bf800043bf000043be800043be000043bd800043bd000043bc800043bc0000",
INIT_30 => X"43c3800043c3000043c2800043c2000043c1800043c1000043c0800043c00000",
INIT_31 => X"43c7800043c7000043c6800043c6000043c5800043c5000043c4800043c40000",
INIT_32 => X"43cb800043cb000043ca800043ca000043c9800043c9000043c8800043c80000",
INIT_33 => X"43cf800043cf000043ce800043ce000043cd800043cd000043cc800043cc0000",
INIT_34 => X"43d3800043d3000043d2800043d2000043d1800043d1000043d0800043d00000",
INIT_35 => X"43d7800043d7000043d6800043d6000043d5800043d5000043d4800043d40000",
INIT_36 => X"43db800043db000043da800043da000043d9800043d9000043d8800043d80000",
INIT_37 => X"43df800043df000043de800043de000043dd800043dd000043dc800043dc0000",
INIT_38 => X"43e3800043e3000043e2800043e2000043e1800043e1000043e0800043e00000",
INIT_39 => X"43e7800043e7000043e6800043e6000043e5800043e5000043e4800043e40000",
INIT_3a => X"43eb800043eb000043ea800043ea000043e9800043e9000043e8800043e80000",
INIT_3b => X"43ef800043ef000043ee800043ee000043ed800043ed000043ec800043ec0000",
INIT_3c => X"43f3800043f3000043f2800043f2000043f1800043f1000043f0800043f00000",
INIT_3d => X"43f7800043f7000043f6800043f6000043f5800043f5000043f4800043f40000",
INIT_3e => X"43fb800043fb000043fa800043fa000043f9800043f9000043f8800043f80000",
INIT_3f => X"43ff800043ff000043fe800043fe000043fd800043fd000043fc800043fc0000",
INIT_40 => X"c3fc8000c3fd0000c3fd8000c3fe0000c3fe8000c3ff0000c3ff8000c4000000",
INIT_41 => X"c3f88000c3f90000c3f98000c3fa0000c3fa8000c3fb0000c3fb8000c3fc0000",
INIT_42 => X"c3f48000c3f50000c3f58000c3f60000c3f68000c3f70000c3f78000c3f80000",
INIT_43 => X"c3f08000c3f10000c3f18000c3f20000c3f28000c3f30000c3f38000c3f40000",
INIT_44 => X"c3ec8000c3ed0000c3ed8000c3ee0000c3ee8000c3ef0000c3ef8000c3f00000",
INIT_45 => X"c3e88000c3e90000c3e98000c3ea0000c3ea8000c3eb0000c3eb8000c3ec0000",
INIT_46 => X"c3e48000c3e50000c3e58000c3e60000c3e68000c3e70000c3e78000c3e80000",
INIT_47 => X"c3e08000c3e10000c3e18000c3e20000c3e28000c3e30000c3e38000c3e40000",
INIT_48 => X"c3dc8000c3dd0000c3dd8000c3de0000c3de8000c3df0000c3df8000c3e00000",
INIT_49 => X"c3d88000c3d90000c3d98000c3da0000c3da8000c3db0000c3db8000c3dc0000",
INIT_4a => X"c3d48000c3d50000c3d58000c3d60000c3d68000c3d70000c3d78000c3d80000",
INIT_4b => X"c3d08000c3d10000c3d18000c3d20000c3d28000c3d30000c3d38000c3d40000",
INIT_4c => X"c3cc8000c3cd0000c3cd8000c3ce0000c3ce8000c3cf0000c3cf8000c3d00000",
INIT_4d => X"c3c88000c3c90000c3c98000c3ca0000c3ca8000c3cb0000c3cb8000c3cc0000",
INIT_4e => X"c3c48000c3c50000c3c58000c3c60000c3c68000c3c70000c3c78000c3c80000",
INIT_4f => X"c3c08000c3c10000c3c18000c3c20000c3c28000c3c30000c3c38000c3c40000",
INIT_50 => X"c3bc8000c3bd0000c3bd8000c3be0000c3be8000c3bf0000c3bf8000c3c00000",
INIT_51 => X"c3b88000c3b90000c3b98000c3ba0000c3ba8000c3bb0000c3bb8000c3bc0000",
INIT_52 => X"c3b48000c3b50000c3b58000c3b60000c3b68000c3b70000c3b78000c3b80000",
INIT_53 => X"c3b08000c3b10000c3b18000c3b20000c3b28000c3b30000c3b38000c3b40000",
INIT_54 => X"c3ac8000c3ad0000c3ad8000c3ae0000c3ae8000c3af0000c3af8000c3b00000",
INIT_55 => X"c3a88000c3a90000c3a98000c3aa0000c3aa8000c3ab0000c3ab8000c3ac0000",
INIT_56 => X"c3a48000c3a50000c3a58000c3a60000c3a68000c3a70000c3a78000c3a80000",
INIT_57 => X"c3a08000c3a10000c3a18000c3a20000c3a28000c3a30000c3a38000c3a40000",
INIT_58 => X"c39c8000c39d0000c39d8000c39e0000c39e8000c39f0000c39f8000c3a00000",
INIT_59 => X"c3988000c3990000c3998000c39a0000c39a8000c39b0000c39b8000c39c0000",
INIT_5a => X"c3948000c3950000c3958000c3960000c3968000c3970000c3978000c3980000",
INIT_5b => X"c3908000c3910000c3918000c3920000c3928000c3930000c3938000c3940000",
INIT_5c => X"c38c8000c38d0000c38d8000c38e0000c38e8000c38f0000c38f8000c3900000",
INIT_5d => X"c3888000c3890000c3898000c38a0000c38a8000c38b0000c38b8000c38c0000",
INIT_5e => X"c3848000c3850000c3858000c3860000c3868000c3870000c3878000c3880000",
INIT_5f => X"c3808000c3810000c3818000c3820000c3828000c3830000c3838000c3840000",
INIT_60 => X"c3790000c37a0000c37b0000c37c0000c37d0000c37e0000c37f0000c3800000",
INIT_61 => X"c3710000c3720000c3730000c3740000c3750000c3760000c3770000c3780000",
INIT_62 => X"c3690000c36a0000c36b0000c36c0000c36d0000c36e0000c36f0000c3700000",
INIT_63 => X"c3610000c3620000c3630000c3640000c3650000c3660000c3670000c3680000",
INIT_64 => X"c3590000c35a0000c35b0000c35c0000c35d0000c35e0000c35f0000c3600000",
INIT_65 => X"c3510000c3520000c3530000c3540000c3550000c3560000c3570000c3580000",
INIT_66 => X"c3490000c34a0000c34b0000c34c0000c34d0000c34e0000c34f0000c3500000",
INIT_67 => X"c3410000c3420000c3430000c3440000c3450000c3460000c3470000c3480000",
INIT_68 => X"c3390000c33a0000c33b0000c33c0000c33d0000c33e0000c33f0000c3400000",
INIT_69 => X"c3310000c3320000c3330000c3340000c3350000c3360000c3370000c3380000",
INIT_6a => X"c3290000c32a0000c32b0000c32c0000c32d0000c32e0000c32f0000c3300000",
INIT_6b => X"c3210000c3220000c3230000c3240000c3250000c3260000c3270000c3280000",
INIT_6c => X"c3190000c31a0000c31b0000c31c0000c31d0000c31e0000c31f0000c3200000",
INIT_6d => X"c3110000c3120000c3130000c3140000c3150000c3160000c3170000c3180000",
INIT_6e => X"c3090000c30a0000c30b0000c30c0000c30d0000c30e0000c30f0000c3100000",
INIT_6f => X"c3010000c3020000c3030000c3040000c3050000c3060000c3070000c3080000",
INIT_70 => X"c2f20000c2f40000c2f60000c2f80000c2fa0000c2fc0000c2fe0000c3000000",
INIT_71 => X"c2e20000c2e40000c2e60000c2e80000c2ea0000c2ec0000c2ee0000c2f00000",
INIT_72 => X"c2d20000c2d40000c2d60000c2d80000c2da0000c2dc0000c2de0000c2e00000",
INIT_73 => X"c2c20000c2c40000c2c60000c2c80000c2ca0000c2cc0000c2ce0000c2d00000",
INIT_74 => X"c2b20000c2b40000c2b60000c2b80000c2ba0000c2bc0000c2be0000c2c00000",
INIT_75 => X"c2a20000c2a40000c2a60000c2a80000c2aa0000c2ac0000c2ae0000c2b00000",
INIT_76 => X"c2920000c2940000c2960000c2980000c29a0000c29c0000c29e0000c2a00000",
INIT_77 => X"c2820000c2840000c2860000c2880000c28a0000c28c0000c28e0000c2900000",
INIT_78 => X"c2640000c2680000c26c0000c2700000c2740000c2780000c27c0000c2800000",
INIT_79 => X"c2440000c2480000c24c0000c2500000c2540000c2580000c25c0000c2600000",
INIT_7a => X"c2240000c2280000c22c0000c2300000c2340000c2380000c23c0000c2400000",
INIT_7b => X"c2040000c2080000c20c0000c2100000c2140000c2180000c21c0000c2200000",
INIT_7c => X"c1c80000c1d00000c1d80000c1e00000c1e80000c1f00000c1f80000c2000000",
INIT_7d => X"c1880000c1900000c1980000c1a00000c1a80000c1b00000c1b80000c1c00000",
INIT_7e => X"c1100000c1200000c1300000c1400000c1500000c1600000c1700000c1800000",
INIT_7f => X"bf800000c0000000c0400000c0800000c0a00000c0c00000c0e00000c1000000"
)
PORT MAP (
DO => o_value,
DOP => open,
ADDR => i_value,
CLK => i_clock,
DI => (others => '0'),
DIP => (others => '0'),
EN => '1',
SSR => i_reset,
WE => '0'
);

end Behavioral;

