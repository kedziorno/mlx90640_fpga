library IEEE;
use IEEE.STD_LOGIC_1164.all;

package colormap_pkg is

type rom_type is array (-128 to 127) of std_logic_vector (23 downto 0);
constant colormap_rom : rom_type := (
x"08003f",
x"08003e",
x"08003e",
x"08003e",
x"09003e",
x"09003e",
x"09003e",
x"09003e",
x"09003e",
x"09003e",
x"09003e",
x"0a003e",
x"0a003e",
x"0a003e",
x"0a003e",
x"0a003e",
x"0a003e",
x"0b003e",
x"0b003e",
x"0b003e",
x"0b003e",
x"0b003e",
x"0b003e",
x"0c003d",
x"0c003d",
x"0c003d",
x"0c003d",
x"0c003d",
x"0c003d",
x"0d003d",
x"0d003d",
x"0d003d",
x"0d003d",
x"0d003c",
x"0e003c",
x"0e003c",
x"0e003c",
x"0e003c",
x"0e003c",
x"0e003c",
x"0f003b",
x"0f003b",
x"0f003b",
x"0f003b",
x"0f003b",
x"10003b",
x"10003b",
x"10003a",
x"10003a",
x"11003a",
x"11003a",
x"11003a",
x"11003a",
x"110039",
x"120039",
x"120039",
x"120039",
x"120039",
x"130038",
x"130038",
x"130038",
x"130038",
x"130038",
x"140037",
x"140037",
x"140037",
x"140037",
x"150036",
x"150036",
x"150036",
x"150036",
x"160036",
x"160035",
x"160035",
x"160035",
x"170035",
x"170034",
x"170034",
x"170034",
x"180034",
x"180033",
x"180033",
x"190033",
x"190033",
x"190032",
x"190032",
x"1a0032",
x"1a0032",
x"1a0031",
x"1a0031",
x"1b0031",
x"1b0030",
x"1b0030",
x"1c0030",
x"1c0030",
x"1c002f",
x"1c002f",
x"1d002f",
x"1d002e",
x"1d002e",
x"1d002e",
x"1e002e",
x"1e002d",
x"1e002d",
x"1f002d",
x"1f002d",
x"1f002c",
x"1f002c",
x"20002c",
x"20002b",
x"20002b",
x"21002b",
x"21002a",
x"21002a",
x"22002a",
x"22002a",
x"220029",
x"220029",
x"230029",
x"230028",
x"230028",
x"240028",
x"240028",
x"240027",
x"250027",
x"250027",
x"250026",
x"250026",
x"260026",
x"260025",
x"260025",
x"270025",
x"270025",
x"270024",
x"280024",
x"280024",
x"280023",
x"280023",
x"290023",
x"290022",
x"290022",
x"2a0022",
x"2a0022",
x"2a0021",
x"2a0021",
x"2b0021",
x"2b0020",
x"2b0020",
x"2c0020",
x"2c001f",
x"2c001f",
x"2d001f",
x"2d001f",
x"2d001e",
x"2d001e",
x"2e001e",
x"2e001d",
x"2e001d",
x"2e001d",
x"2f001d",
x"2f001c",
x"2f001c",
x"30001c",
x"30001c",
x"30001b",
x"30001b",
x"31001b",
x"31001a",
x"31001a",
x"32001a",
x"32001a",
x"320019",
x"320019",
x"330019",
x"330019",
x"330018",
x"330018",
x"340018",
x"340017",
x"340017",
x"340017",
x"350017",
x"350016",
x"350016",
x"350016",
x"360016",
x"360015",
x"360015",
x"360015",
x"360015",
x"370014",
x"370014",
x"370014",
x"370014",
x"380013",
x"380013",
x"380013",
x"380013",
x"380013",
x"390012",
x"390012",
x"390012",
x"390012",
x"390011",
x"3a0011",
x"3a0011",
x"3a0011",
x"3a0011",
x"3a0010",
x"3a0010",
x"3b0010",
x"3b0010",
x"3b000f",
x"3b000f",
x"3b000f",
x"3b000f",
x"3b000f",
x"3c000e",
x"3c000e",
x"3c000e",
x"3c000e",
x"3c000e",
x"3c000e",
x"3c000d",
x"3d000d",
x"3d000d",
x"3d000d",
x"3d000d",
x"3d000c",
x"3d000c",
x"3d000c",
x"3d000c",
x"3d000c",
x"3d000c",
x"3e000b",
x"3e000b",
x"3e000b",
x"3e000b",
x"3e000b",
x"3e000b",
x"3e000a",
x"3e000a",
x"3e000a",
x"3e000a",
x"3e000a",
x"3e000a",
x"3e0009",
x"3e0009",
x"3e0009",
x"3e0009",
x"3e0009",
x"3e0009",
x"3e0009",
x"3e0008",
x"3e0008",
x"3e0008"
);

end colormap_pkg;

package body colormap_pkg is
 
end colormap_pkg;
