library IEEE;
use IEEE.STD_LOGIC_1164.all;

package p_package1_constants is


end p_package1_constants;

package body p_package1_constants is


end p_package1_constants;
