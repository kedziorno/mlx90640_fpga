----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:08:59 01/24/2023 
-- Design Name: 
-- Module Name:    ExtractVDDParameters - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

--    RAMB16     : In order to incorporate this function into the design,
--     VHDL      : the following instance declaration needs to be placed
--   instance    : in the architecture body of the design code.  The
--  declaration  : (RAMB16_inst) and/or the port declarations
--     code      : after the "=>" assignment maybe changed to properly
--               : reference and connect this function to the design.
--               : All inputs and outputs must be connected.
--    Library    : In addition to adding the instance declaration, a use
--  declaration  : statement for the UNISIM.vcomponents library needs to be
--      for      : added before the entity declaration.  This library
--    Xilinx     : contains the component declarations for all Xilinx
--   primitives  : primitives and points to the models that will be used
--               : for simulation.
--  Copy the following two statements and paste them before the
--  Entity declaration, unless they already exist.
----  <-----Cut code below this line and paste into the architecture body---->
--
--   -- RAMB16: 16k+2k Parity Parameterizable BlockRAM
--   --         Virtex-4
--   -- Xilinx HDL Language Template, version 14.7
--
--   RAMB16_inst : RAMB16
--   generic map (
--      DOA_REG => 0, -- Optional output registers on the A port (0 or 1)
--      DOB_REG => 0, -- Optional output registers on the B port (0 or 1)
--      INIT_A => X"000000000", --  Initial values on A output port
--      INIT_B => X"000000000", --  Initial values on B output port
--      INVERT_CLK_DOA_REG => FALSE, -- Invert clock on A port output registers (TRUE or FALSE)
--      INVERT_CLK_DOB_REG => FALSE, -- Invert clock on B port output registers (TRUE or FALSE)
--      RAM_EXTENSION_A => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--      RAM_EXTENSION_B => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
--      READ_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36 
--      READ_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36 
--      SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
--                                    -- "GENERATE_X_ONLY" or "NONE" 
--      SRVAL_A => X"000000000", --  Port A output value upon SSR assertion
--      SRVAL_B => X"000000000", --  Port B output value upon SSR assertion
--      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
--      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
--      WRITE_WIDTH_A => 0, -- Valid values are 1,2,4,9,18 or 36
--      WRITE_WIDTH_B => 0, -- Valid values are 1,2,4,9,18 or 36 
--      -- The following INIT_xx declarations specify the initial contents of the RAM
--      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
--      -- The next set of INITP_xx are for the parity bits
--      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
--   port map (
--      CASCADEOUTA => CASCADEOUTA, -- 1-bit cascade output
--      CASCADEOUTB => CASCADEOUTB, -- 1-bit cascade output
--      DOA => DOA,      -- 32-bit A port Data Output
--      DOB => DOB,      -- 32-bit B port Data Output
--      DOPA => DOPA,    -- 4-bit  A port Parity Output
--      DOPB => DOPB,    -- 4-bit  B port Parity Output
--      ADDRA => ADDRA,  -- 15-bit A port Address Input
--      ADDRB => ADDRB,  -- 15-bit B port Address Input
--      CASCADEINA => CASCADEINA, -- 1-bit cascade A input
--      CASCADEINB => CASCADEINB, -- 1-bit cascade B input
--      CLKA => CLKA,    -- Port A Clock
--      CLKB => CLKB,    -- Port B Clock
--      DIA => DIA,      -- 32-bit A port Data Input
--      DIB => DIB,      -- 32-bit B port Data Input
--      DIPA => DIPA,    -- 4-bit  A port parity Input
--      DIPB => DIPB,    -- 4-bit  B port parity Input
--      ENA => ENA,      -- 1-bit  A port Enable Input
--      ENB => ENB,      -- 1-bit  B port Enable Input
--      REGCEA => REGCEA, -- 1-bit A port register enable input
--      REGCEB => REGCEB, -- 1-bit B port register enable input
--      SSRA => SSRA,    -- 1-bit  A port Synchronous Set/Reset Input
--      SSRB => SSRB,    -- 1-bit  B port Synchronous Set/Reset Input
--      WEA => WEA,      -- 4-bit  A port Write Enable Input
--      WEB => WEB       -- 4-bit  B port Write Enable Input
--   );
--
--   -- End of RAMB16_inst instantiation

entity ExtractVDDParameters is
port (
i_clock : IN  std_logic;
i_reset : IN  std_logic;
i_run : in std_logic;
i2c_mem_ena : out STD_LOGIC;
i2c_mem_addra : out STD_LOGIC_VECTOR(11 DOWNTO 0);
i2c_mem_douta : in STD_LOGIC_VECTOR(7 DOWNTO 0);
o_kvdd : OUT  std_logic_vector (31 downto 0);
o_vdd25 : OUT  std_logic_vector (31 downto 0);
o_rdy : out std_logic
);
end ExtractVDDParameters;

architecture Behavioral of ExtractVDDParameters is

--component RAMB16 is
--  generic (
--    DOA_REG : integer := 0 ;
--    DOB_REG : integer := 0 ;
--    INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INIT_A : bit_vector := X"000000000";
--    INIT_B : bit_vector := X"000000000";
--    INIT_FILE : string := "NONE";
--    INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
--    INVERT_CLK_DOA_REG : boolean := false;
--    INVERT_CLK_DOB_REG : boolean := false;
--    RAM_EXTENSION_A : string := "NONE";
--    RAM_EXTENSION_B : string := "NONE";
--    READ_WIDTH_A : integer := 18;
--    READ_WIDTH_B : integer := 18;
--    SIM_COLLISION_CHECK : string := "ALL";
--    SRVAL_A  : bit_vector := X"000000000";
--    SRVAL_B  : bit_vector := X"000000000";
--    WRITE_MODE_A : string := "WRITE_FIRST";
--    WRITE_MODE_B : string := "WRITE_FIRST";
--    WRITE_WIDTH_A : integer := 0;
--    WRITE_WIDTH_B : integer := 0
--  );
--  port(
--    CASCADEOUTA  : out  std_ulogic;
--    CASCADEOUTB  : out  std_ulogic;
--    DOA          : out std_logic_vector (31 downto 0);
--    DOB          : out std_logic_vector (31 downto 0);
--    DOPA         : out std_logic_vector (3 downto 0);
--    DOPB         : out std_logic_vector (3 downto 0);
--    ADDRA        : in  std_logic_vector (14 downto 0);
--    ADDRB        : in  std_logic_vector (14 downto 0);
--    CASCADEINA   : in  std_ulogic := '0';
--    CASCADEINB   : in  std_ulogic := '0';
--    CLKA         : in  std_ulogic;
--    CLKB         : in  std_ulogic;
--    DIA          : in  std_logic_vector (31 downto 0) := (others => '0');
--    DIB          : in  std_logic_vector (31 downto 0) := (others => '0');
--    DIPA         : in  std_logic_vector (3 downto 0) := (others => '0');
--    DIPB         : in  std_logic_vector (3 downto 0) := (others => '0');
--    ENA          : in  std_ulogic := '0';
--    ENB          : in  std_ulogic := '0';
--    REGCEA       : in  std_ulogic := '0';
--    REGCEB       : in  std_ulogic := '0';
--    SSRA         : in  std_ulogic := '0';
--    SSRB         : in  std_ulogic := '0';
--    WEA          : in  std_logic_vector (3 downto 0) := (others => '0');
--    WEB          : in  std_logic_vector (3 downto 0) := (others => '0')
--  );
--end component RAMB16;

signal odata_kvdd : std_logic_vector (31 downto 0);
signal odata_vdd25 : std_logic_vector (31 downto 0);
--signal address_kvdd : std_logic_vector (14 downto 0);
--signal address_vdd25 : std_logic_vector (14 downto 0);
signal address_kvdd : std_logic_vector (8 downto 0);
signal address_vdd25 : std_logic_vector (8 downto 0);

begin

p0 : process (i_clock) is
	variable ee2433 : std_logic_vector (15 downto 0);
	type states is (idle,s1,s2,s3,s4,s5,s6,s7,ending);
	variable state : states;
begin
	if (rising_edge (i_clock)) then
		if (i_reset = '1') then
			state := idle;
			i2c_mem_ena <= '0';
			o_rdy <= '0';
		else
			case (state) is
				when idle =>
					if (i_run = '1') then
						state := s1;
						i2c_mem_ena <= '1';
					else
						state := idle;
						i2c_mem_ena <= '0';
					end if;
				when s1 => state := s2;
					i2c_mem_addra <= std_logic_vector (to_unsigned (51*2+0, 12)); -- 2433 MSB kvdd
				when s2 => state := s3;
					i2c_mem_addra <= std_logic_vector (to_unsigned (51*2+1, 12)); -- 2433 LSB vdd25
				when s3 => state := s4;
					ee2433 (15 downto 8) := i2c_mem_douta;
				when s4 => state := s5;
					ee2433 (7 downto 0) := i2c_mem_douta;
				when s5 => state := s6;
					address_kvdd  <= "0"&ee2433 (15 downto 8);
					address_vdd25 <= "1"&ee2433 (7 downto 0);
				when s6 => state := s7;
				when s7 => state := ending;
--					o_kvdd <= odata_kvdd (19 downto 0)&x"000";
--					o_vdd25 <= odata_vdd25 (19 downto 0)&x"000";
					o_kvdd <= odata_kvdd;
					o_vdd25 <= odata_vdd25;
				when ending => state := idle;
					o_rdy <= '1';
			end case;
		end if;
	end if;
end process p0;

inst_mem_kvdd_vdd25 : RAMB16_S36_S36 -- XXX on xc4vsx35 syn not work (RAMB16)
generic map (
INIT_A => X"000000000", -- Value of output RAM registers on Port A at startup
INIT_B => X"000000000", -- Value of output RAM registers on Port B at startup
SRVAL_A => X"000000000", -- Port A output value upon SSR assertion
SRVAL_B => X"000000000", -- Port B output value upon SSR assertion
WRITE_MODE_A => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
WRITE_MODE_B => "WRITE_FIRST", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
SIM_COLLISION_CHECK => "NONE", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"-- The following INIT_xx declarations specify the intial contents of the RAM

INIT_00 => X"4360000043400000432000004300000042c00000428000004200000022000000", -- 43000000
INIT_01 => X"43f0000043e0000043d0000043c0000043b0000043a000004390000043800000", -- 43b00000
INIT_02 => X"4438000044300000442800004420000044180000441000004408000044000000",
INIT_03 => X"4478000044700000446800004460000044580000445000004448000044400000",
INIT_04 => X"449c0000449800004494000044900000448c0000448800004484000044800000",
INIT_05 => X"44bc000044b8000044b4000044b0000044ac000044a8000044a4000044a00000",
INIT_06 => X"44dc000044d8000044d4000044d0000044cc000044c8000044c4000044c00000",
INIT_07 => X"44fc000044f8000044f4000044f0000044ec000044e8000044e4000044e00000",
INIT_08 => X"450e0000450c0000450a00004508000045060000450400004502000045000000",
INIT_09 => X"451e0000451c0000451a00004518000045160000451400004512000045100000",
INIT_0a => X"452e0000452c0000452a00004528000045260000452400004522000045200000",
INIT_0b => X"453e0000453c0000453a00004538000045360000453400004532000045300000",
INIT_0c => X"454e0000454c0000454a00004548000045460000454400004542000045400000",
INIT_0d => X"455e0000455c0000455a00004558000045560000455400004552000045500000",
INIT_0e => X"456e0000456c0000456a00004568000045660000456400004562000045600000",
INIT_0f => X"457e0000457c0000457a00004578000045760000457400004572000045700000",
INIT_10 => X"c5720000c5740000c5760000c5780000c57a0000c57c0000c57e0000c5800000",
INIT_11 => X"c5620000c5640000c5660000c5680000c56a0000c56c0000c56e0000c5700000",
INIT_12 => X"c5520000c5540000c5560000c5580000c55a0000c55c0000c55e0000c5600000",
INIT_13 => X"c5420000c5440000c5460000c5480000c54a0000c54c0000c54e0000c5500000",--
INIT_14 => X"c5320000c5340000c5360000c5380000c53a0000c53c0000c53e0000c5400000",
INIT_15 => X"c5220000c5240000c5260000c5280000c52a0000c52c0000c52e0000c5300000",
INIT_16 => X"c5120000c5140000c5160000c5180000c51a0000c51c0000c51e0000c5200000",
INIT_17 => X"c5020000c5040000c5060000c5080000c50a0000c50c0000c50e0000c5100000",
INIT_18 => X"c4e40000c4e80000c4ec0000c4f00000c4f40000c4f80000c4fc0000c5000000",
INIT_19 => X"c4c40000c4c80000c4cc0000c4d00000c4d40000c4d80000c4dc0000c4e00000",
INIT_1a => X"c4a40000c4a80000c4ac0000c4b00000c4b40000c4b80000c4bc0000c4c00000",
INIT_1b => X"c4840000c4880000c48c0000c4900000c4940000c4980000c49c0000c4a00000",
INIT_1c => X"c4480000c4500000c4580000c4600000c4680000c4700000c4780000c4800000",
INIT_1d => X"c4080000c4100000c4180000c4200000c4280000c4300000c4380000c4400000",
INIT_1e => X"c3900000c3a00000c3b00000c3c00000c3d00000c3e00000c3f00000c4000000",
INIT_1f => X"c2000000c2800000c2c00000c3000000c3200000c3400000c3600000c3800000",

INIT_20 => X"c67c8000c67d0000c67d8000c67e0000c67e8000c67f0000c67f8000c6800000",
INIT_21 => X"c6788000c6790000c6798000c67a0000c67a8000c67b0000c67b8000c67c0000",
INIT_22 => X"c6748000c6750000c6758000c6760000c6768000c6770000c6778000c6780000",
INIT_23 => X"c6708000c6710000c6718000c6720000c6728000c6730000c6738000c6740000",
INIT_24 => X"c66c8000c66d0000c66d8000c66e0000c66e8000c66f0000c66f8000c6700000",
INIT_25 => X"c6688000c6690000c6698000c66a0000c66a8000c66b0000c66b8000c66c0000",
INIT_26 => X"c6648000c6650000c6658000c6660000c6668000c6670000c6678000c6680000",
INIT_27 => X"c6608000c6610000c6618000c6620000c6628000c6630000c6638000c6640000",
INIT_28 => X"c65c8000c65d0000c65d8000c65e0000c65e8000c65f0000c65f8000c6600000",
INIT_29 => X"c6588000c6590000c6598000c65a0000c65a8000c65b0000c65b8000c65c0000",
INIT_2a => X"c6548000c6550000c6558000c6560000c6568000c6570000c6578000c6580000",
INIT_2b => X"c6508000c6510000c6518000c6520000c6528000c6530000c6538000c6540000",
INIT_2c => X"c64c8000c64d0000c64d8000c64e0000c64e8000c64f0000c64f8000c6500000",
INIT_2d => X"c6488000c6490000c6498000c64a0000c64a8000c64b0000c64b8000c64c0000", -- c64c0000
INIT_2e => X"c6448000c6450000c6458000c6460000c6468000c6470000c6478000c6480000",
INIT_2f => X"c6408000c6410000c6418000c6420000c6428000c6430000c6438000c6440000",
INIT_30 => X"c63c8000c63d0000c63d8000c63e0000c63e8000c63f0000c63f8000c6400000",
INIT_31 => X"c6388000c6390000c6398000c63a0000c63a8000c63b0000c63b8000c63c0000",
INIT_32 => X"c6348000c6350000c6358000c6360000c6368000c6370000c6378000c6380000",
INIT_33 => X"c6308000c6310000c6318000c6320000c6328000c6330000c6338000c6340000",
INIT_34 => X"c62c8000c62d0000c62d8000c62e0000c62e8000c62f0000c62f8000c6300000",
INIT_35 => X"c6288000c6290000c6298000c62a0000c62a8000c62b0000c62b8000c62c0000",
INIT_36 => X"c6248000c6250000c6258000c6260000c6268000c6270000c6278000c6280000",
INIT_37 => X"c6208000c6210000c6218000c6220000c6228000c6230000c6238000c6240000",
INIT_38 => X"c61c8000c61d0000c61d8000c61e0000c61e8000c61f0000c61f8000c6200000",
INIT_39 => X"c6188000c6190000c6198000c61a0000c61a8000c61b0000c61b8000c61c0000",
INIT_3a => X"c6148000c6150000c6158000c6160000c6168000c6170000c6178000c6180000",
INIT_3b => X"c6108000c6110000c6118000c6120000c6128000c6130000c6138000c6140000",
INIT_3c => X"c60c8000c60d0000c60d8000c60e0000c60e8000c60f0000c60f8000c6100000",
INIT_3d => X"c6088000c6090000c6098000c60a0000c60a8000c60b0000c60b8000c60c0000",
INIT_3e => X"c6048000c6050000c6058000c6060000c6068000c6070000c6078000c6080000",
INIT_3f => X"c6008000c6010000c6018000c6020000c6028000c6030000c6038000c6040000"
)
port map (
DOA => odata_kvdd, -- 1-bit Data Output
DOPA => open, -- 1-bit Data Output
ADDRA => address_kvdd, -- 14-bit Address Input
CLKA => i_clock, -- Clock
DIA => (others => '0'), -- 1-bit Data Input
DIPA => (others => '0'), -- 1-bit Data Input
ENA => '1', -- RAM Enable Input
SSRA => i_reset, -- Synchronous Set/Reset Input
WEA => '0', -- Write Enable Input,

DOB => odata_vdd25, -- 1-bit Data Output
DOPB => open, -- 1-bit Data Output
ADDRB => address_vdd25, -- 14-bit Address Input
CLKB => i_clock, -- Clock
DIB => (others => '0'), -- 1-bit Data Input
DIPB => (others => '0'), -- 1-bit Data Input
ENB => '1', -- RAM Enable Input
SSRB => i_reset, -- Synchronous Set/Reset Input
WEB => '0' -- Write Enable Input,
);

end Behavioral;
